magic
tech scmos
timestamp 1636179762
<< ab >>
rect 0 5 87 77
rect 91 39 218 77
rect 91 30 128 39
rect 131 30 218 39
rect 91 26 218 30
rect 91 24 129 26
rect 131 24 218 26
rect 91 5 218 24
rect 220 39 347 77
rect 220 30 307 39
rect 310 30 347 39
rect 220 26 347 30
rect 220 24 307 26
rect 309 24 347 26
rect 220 5 347 24
rect 351 5 525 77
rect 529 39 751 77
rect 529 30 566 39
rect 569 30 751 39
rect 529 26 751 30
rect 529 24 567 26
rect 569 24 751 26
rect 529 5 751 24
<< nwell >>
rect 0 37 751 82
<< pwell >>
rect 0 0 751 37
<< poly >>
rect 10 71 12 75
rect 20 71 22 75
rect 30 71 32 75
rect 48 68 50 73
rect 55 68 57 73
rect 78 71 80 75
rect 98 71 100 75
rect 105 71 107 75
rect 65 59 67 64
rect 139 71 141 75
rect 149 71 151 75
rect 159 71 161 75
rect 118 62 120 66
rect 65 43 67 46
rect 10 40 12 43
rect 20 40 22 43
rect 30 40 32 43
rect 48 40 50 43
rect 55 40 57 43
rect 65 41 74 43
rect 8 38 14 40
rect 8 36 10 38
rect 12 36 14 38
rect 8 34 14 36
rect 18 38 24 40
rect 18 36 20 38
rect 22 36 24 38
rect 18 34 24 36
rect 28 38 50 40
rect 28 36 30 38
rect 32 36 37 38
rect 39 36 50 38
rect 28 34 50 36
rect 54 38 60 40
rect 54 36 56 38
rect 58 36 60 38
rect 54 34 60 36
rect 10 25 12 34
rect 21 31 23 34
rect 28 31 30 34
rect 48 31 50 34
rect 58 31 60 34
rect 68 39 70 41
rect 72 39 74 41
rect 68 37 74 39
rect 68 24 70 37
rect 78 33 80 46
rect 98 40 100 53
rect 105 48 107 53
rect 104 46 110 48
rect 104 44 106 46
rect 108 44 110 46
rect 104 42 110 44
rect 94 38 100 40
rect 94 36 96 38
rect 98 36 100 38
rect 94 34 100 36
rect 74 31 80 33
rect 74 29 76 31
rect 78 29 80 31
rect 74 27 80 29
rect 78 24 80 27
rect 98 26 100 34
rect 108 26 110 42
rect 118 41 120 50
rect 177 68 179 73
rect 184 68 186 73
rect 207 71 209 75
rect 229 71 231 75
rect 194 59 196 64
rect 252 68 254 73
rect 259 68 261 73
rect 277 71 279 75
rect 287 71 289 75
rect 297 71 299 75
rect 242 59 244 64
rect 194 43 196 46
rect 114 39 120 41
rect 139 40 141 43
rect 149 40 151 43
rect 159 40 161 43
rect 177 40 179 43
rect 184 40 186 43
rect 194 41 203 43
rect 114 37 116 39
rect 118 37 120 39
rect 114 35 120 37
rect 118 26 120 35
rect 137 38 143 40
rect 137 36 139 38
rect 141 36 143 38
rect 137 34 143 36
rect 147 38 153 40
rect 147 36 149 38
rect 151 36 153 38
rect 147 34 153 36
rect 157 38 179 40
rect 157 36 159 38
rect 161 36 166 38
rect 168 36 179 38
rect 157 34 179 36
rect 183 38 189 40
rect 183 36 185 38
rect 187 36 189 38
rect 183 34 189 36
rect 48 12 50 17
rect 58 12 60 17
rect 10 7 12 11
rect 21 7 23 11
rect 28 7 30 11
rect 68 9 70 14
rect 139 25 141 34
rect 150 31 152 34
rect 157 31 159 34
rect 177 31 179 34
rect 187 31 189 34
rect 197 39 199 41
rect 201 39 203 41
rect 197 37 203 39
rect 98 16 100 20
rect 108 16 110 20
rect 118 16 120 20
rect 78 7 80 11
rect 197 24 199 37
rect 207 33 209 46
rect 203 31 209 33
rect 203 29 205 31
rect 207 29 209 31
rect 203 27 209 29
rect 207 24 209 27
rect 229 33 231 46
rect 242 43 244 46
rect 331 71 333 75
rect 338 71 340 75
rect 358 71 360 75
rect 318 62 320 66
rect 235 41 244 43
rect 235 39 237 41
rect 239 39 241 41
rect 252 40 254 43
rect 259 40 261 43
rect 277 40 279 43
rect 287 40 289 43
rect 297 40 299 43
rect 318 41 320 50
rect 331 48 333 53
rect 328 46 334 48
rect 328 44 330 46
rect 332 44 334 46
rect 328 42 334 44
rect 235 37 241 39
rect 229 31 235 33
rect 229 29 231 31
rect 233 29 235 31
rect 229 27 235 29
rect 229 24 231 27
rect 239 24 241 37
rect 249 38 255 40
rect 249 36 251 38
rect 253 36 255 38
rect 249 34 255 36
rect 259 38 281 40
rect 259 36 270 38
rect 272 36 277 38
rect 279 36 281 38
rect 259 34 281 36
rect 285 38 291 40
rect 285 36 287 38
rect 289 36 291 38
rect 285 34 291 36
rect 295 38 301 40
rect 295 36 297 38
rect 299 36 301 38
rect 295 34 301 36
rect 318 39 324 41
rect 318 37 320 39
rect 322 37 324 39
rect 318 35 324 37
rect 249 31 251 34
rect 259 31 261 34
rect 279 31 281 34
rect 286 31 288 34
rect 177 12 179 17
rect 187 12 189 17
rect 139 7 141 11
rect 150 7 152 11
rect 157 7 159 11
rect 197 9 199 14
rect 207 7 209 11
rect 229 7 231 11
rect 239 9 241 14
rect 249 12 251 17
rect 259 12 261 17
rect 297 25 299 34
rect 318 26 320 35
rect 328 26 330 42
rect 338 40 340 53
rect 381 68 383 73
rect 388 68 390 73
rect 406 71 408 75
rect 416 71 418 75
rect 426 71 428 75
rect 448 71 450 75
rect 458 71 460 75
rect 468 71 470 75
rect 371 59 373 64
rect 338 38 344 40
rect 338 36 340 38
rect 342 36 344 38
rect 338 34 344 36
rect 338 26 340 34
rect 358 33 360 46
rect 371 43 373 46
rect 486 68 488 73
rect 493 68 495 73
rect 516 71 518 75
rect 536 71 538 75
rect 543 71 545 75
rect 503 59 505 64
rect 577 71 579 75
rect 587 71 589 75
rect 597 71 599 75
rect 556 62 558 66
rect 503 43 505 46
rect 364 41 373 43
rect 364 39 366 41
rect 368 39 370 41
rect 381 40 383 43
rect 388 40 390 43
rect 406 40 408 43
rect 416 40 418 43
rect 426 40 428 43
rect 448 40 450 43
rect 458 40 460 43
rect 468 40 470 43
rect 486 40 488 43
rect 493 40 495 43
rect 503 41 512 43
rect 364 37 370 39
rect 358 31 364 33
rect 358 29 360 31
rect 362 29 364 31
rect 358 27 364 29
rect 358 24 360 27
rect 368 24 370 37
rect 378 38 384 40
rect 378 36 380 38
rect 382 36 384 38
rect 378 34 384 36
rect 388 38 410 40
rect 388 36 399 38
rect 401 36 406 38
rect 408 36 410 38
rect 388 34 410 36
rect 414 38 420 40
rect 414 36 416 38
rect 418 36 420 38
rect 414 34 420 36
rect 424 38 430 40
rect 424 36 426 38
rect 428 36 430 38
rect 424 34 430 36
rect 446 38 452 40
rect 446 36 448 38
rect 450 36 452 38
rect 446 34 452 36
rect 456 38 462 40
rect 456 36 458 38
rect 460 36 462 38
rect 456 34 462 36
rect 466 38 488 40
rect 466 36 468 38
rect 470 36 475 38
rect 477 36 488 38
rect 466 34 488 36
rect 492 38 498 40
rect 492 36 494 38
rect 496 36 498 38
rect 492 34 498 36
rect 378 31 380 34
rect 388 31 390 34
rect 408 31 410 34
rect 415 31 417 34
rect 318 16 320 20
rect 328 16 330 20
rect 338 16 340 20
rect 279 7 281 11
rect 286 7 288 11
rect 297 7 299 11
rect 358 7 360 11
rect 368 9 370 14
rect 378 12 380 17
rect 388 12 390 17
rect 426 25 428 34
rect 448 25 450 34
rect 459 31 461 34
rect 466 31 468 34
rect 486 31 488 34
rect 496 31 498 34
rect 506 39 508 41
rect 510 39 512 41
rect 506 37 512 39
rect 506 24 508 37
rect 516 33 518 46
rect 536 40 538 53
rect 543 48 545 53
rect 542 46 548 48
rect 542 44 544 46
rect 546 44 548 46
rect 542 42 548 44
rect 532 38 538 40
rect 532 36 534 38
rect 536 36 538 38
rect 532 34 538 36
rect 512 31 518 33
rect 512 29 514 31
rect 516 29 518 31
rect 512 27 518 29
rect 516 24 518 27
rect 536 26 538 34
rect 546 26 548 42
rect 556 41 558 50
rect 615 68 617 73
rect 622 68 624 73
rect 645 71 647 75
rect 669 71 671 75
rect 679 71 681 75
rect 689 71 691 75
rect 632 59 634 64
rect 632 43 634 46
rect 552 39 558 41
rect 577 40 579 43
rect 587 40 589 43
rect 597 40 599 43
rect 615 40 617 43
rect 622 40 624 43
rect 632 41 641 43
rect 552 37 554 39
rect 556 37 558 39
rect 552 35 558 37
rect 556 26 558 35
rect 575 38 581 40
rect 575 36 577 38
rect 579 36 581 38
rect 575 34 581 36
rect 585 38 591 40
rect 585 36 587 38
rect 589 36 591 38
rect 585 34 591 36
rect 595 38 617 40
rect 595 36 597 38
rect 599 36 604 38
rect 606 36 617 38
rect 595 34 617 36
rect 621 38 627 40
rect 621 36 623 38
rect 625 36 627 38
rect 621 34 627 36
rect 486 12 488 17
rect 496 12 498 17
rect 408 7 410 11
rect 415 7 417 11
rect 426 7 428 11
rect 448 7 450 11
rect 459 7 461 11
rect 466 7 468 11
rect 506 9 508 14
rect 577 25 579 34
rect 588 31 590 34
rect 595 31 597 34
rect 615 31 617 34
rect 625 31 627 34
rect 635 39 637 41
rect 639 39 641 41
rect 635 37 641 39
rect 536 16 538 20
rect 546 16 548 20
rect 556 16 558 20
rect 516 7 518 11
rect 635 24 637 37
rect 645 33 647 46
rect 707 68 709 73
rect 714 68 716 73
rect 737 71 739 75
rect 724 59 726 64
rect 724 43 726 46
rect 669 40 671 43
rect 679 40 681 43
rect 689 40 691 43
rect 707 40 709 43
rect 714 40 716 43
rect 724 41 733 43
rect 667 38 673 40
rect 667 36 669 38
rect 671 36 673 38
rect 667 34 673 36
rect 677 38 683 40
rect 677 36 679 38
rect 681 36 683 38
rect 677 34 683 36
rect 687 38 709 40
rect 687 36 689 38
rect 691 36 696 38
rect 698 36 709 38
rect 687 34 709 36
rect 713 38 719 40
rect 713 36 715 38
rect 717 36 719 38
rect 713 34 719 36
rect 641 31 647 33
rect 641 29 643 31
rect 645 29 647 31
rect 641 27 647 29
rect 645 24 647 27
rect 669 25 671 34
rect 680 31 682 34
rect 687 31 689 34
rect 707 31 709 34
rect 717 31 719 34
rect 727 39 729 41
rect 731 39 733 41
rect 727 37 733 39
rect 615 12 617 17
rect 625 12 627 17
rect 577 7 579 11
rect 588 7 590 11
rect 595 7 597 11
rect 635 9 637 14
rect 727 24 729 37
rect 737 33 739 46
rect 733 31 739 33
rect 733 29 735 31
rect 737 29 739 31
rect 733 27 739 29
rect 737 24 739 27
rect 707 12 709 17
rect 717 12 719 17
rect 645 7 647 11
rect 669 7 671 11
rect 680 7 682 11
rect 687 7 689 11
rect 727 9 729 14
rect 737 7 739 11
<< ndif >>
rect 14 25 21 31
rect 3 22 10 25
rect 3 20 5 22
rect 7 20 10 22
rect 3 18 10 20
rect 5 11 10 18
rect 12 15 21 25
rect 12 13 16 15
rect 18 13 21 15
rect 12 11 21 13
rect 23 11 28 31
rect 30 24 35 31
rect 41 29 48 31
rect 41 27 43 29
rect 45 27 48 29
rect 30 22 37 24
rect 30 20 33 22
rect 35 20 37 22
rect 30 18 37 20
rect 41 22 48 27
rect 41 20 43 22
rect 45 20 48 22
rect 30 11 35 18
rect 41 17 48 20
rect 50 29 58 31
rect 50 27 53 29
rect 55 27 58 29
rect 50 17 58 27
rect 60 24 65 31
rect 91 24 98 26
rect 60 21 68 24
rect 60 19 63 21
rect 65 19 68 21
rect 60 17 68 19
rect 63 14 68 17
rect 70 18 78 24
rect 70 16 73 18
rect 75 16 78 18
rect 70 14 78 16
rect 73 11 78 14
rect 80 22 87 24
rect 80 20 83 22
rect 85 20 87 22
rect 91 22 93 24
rect 95 22 98 24
rect 91 20 98 22
rect 100 24 108 26
rect 100 22 103 24
rect 105 22 108 24
rect 100 20 108 22
rect 110 24 118 26
rect 110 22 113 24
rect 115 22 118 24
rect 110 20 118 22
rect 120 24 127 26
rect 143 25 150 31
rect 120 22 123 24
rect 125 22 127 24
rect 120 20 127 22
rect 132 22 139 25
rect 132 20 134 22
rect 136 20 139 22
rect 80 18 87 20
rect 80 11 85 18
rect 132 18 139 20
rect 134 11 139 18
rect 141 15 150 25
rect 141 13 145 15
rect 147 13 150 15
rect 141 11 150 13
rect 152 11 157 31
rect 159 24 164 31
rect 170 29 177 31
rect 170 27 172 29
rect 174 27 177 29
rect 159 22 166 24
rect 159 20 162 22
rect 164 20 166 22
rect 159 18 166 20
rect 170 22 177 27
rect 170 20 172 22
rect 174 20 177 22
rect 159 11 164 18
rect 170 17 177 20
rect 179 29 187 31
rect 179 27 182 29
rect 184 27 187 29
rect 179 17 187 27
rect 189 24 194 31
rect 244 24 249 31
rect 189 21 197 24
rect 189 19 192 21
rect 194 19 197 21
rect 189 17 197 19
rect 192 14 197 17
rect 199 18 207 24
rect 199 16 202 18
rect 204 16 207 18
rect 199 14 207 16
rect 202 11 207 14
rect 209 22 216 24
rect 209 20 212 22
rect 214 20 216 22
rect 209 18 216 20
rect 222 22 229 24
rect 222 20 224 22
rect 226 20 229 22
rect 222 18 229 20
rect 209 11 214 18
rect 224 11 229 18
rect 231 18 239 24
rect 231 16 234 18
rect 236 16 239 18
rect 231 14 239 16
rect 241 21 249 24
rect 241 19 244 21
rect 246 19 249 21
rect 241 17 249 19
rect 251 29 259 31
rect 251 27 254 29
rect 256 27 259 29
rect 251 17 259 27
rect 261 29 268 31
rect 261 27 264 29
rect 266 27 268 29
rect 261 22 268 27
rect 274 24 279 31
rect 261 20 264 22
rect 266 20 268 22
rect 261 17 268 20
rect 272 22 279 24
rect 272 20 274 22
rect 276 20 279 22
rect 272 18 279 20
rect 241 14 246 17
rect 231 11 236 14
rect 274 11 279 18
rect 281 11 286 31
rect 288 25 295 31
rect 288 15 297 25
rect 288 13 291 15
rect 293 13 297 15
rect 288 11 297 13
rect 299 22 306 25
rect 299 20 302 22
rect 304 20 306 22
rect 311 24 318 26
rect 311 22 313 24
rect 315 22 318 24
rect 311 20 318 22
rect 320 24 328 26
rect 320 22 323 24
rect 325 22 328 24
rect 320 20 328 22
rect 330 24 338 26
rect 330 22 333 24
rect 335 22 338 24
rect 330 20 338 22
rect 340 24 347 26
rect 373 24 378 31
rect 340 22 343 24
rect 345 22 347 24
rect 340 20 347 22
rect 351 22 358 24
rect 351 20 353 22
rect 355 20 358 22
rect 299 18 306 20
rect 299 11 304 18
rect 351 18 358 20
rect 353 11 358 18
rect 360 18 368 24
rect 360 16 363 18
rect 365 16 368 18
rect 360 14 368 16
rect 370 21 378 24
rect 370 19 373 21
rect 375 19 378 21
rect 370 17 378 19
rect 380 29 388 31
rect 380 27 383 29
rect 385 27 388 29
rect 380 17 388 27
rect 390 29 397 31
rect 390 27 393 29
rect 395 27 397 29
rect 390 22 397 27
rect 403 24 408 31
rect 390 20 393 22
rect 395 20 397 22
rect 390 17 397 20
rect 401 22 408 24
rect 401 20 403 22
rect 405 20 408 22
rect 401 18 408 20
rect 370 14 375 17
rect 360 11 365 14
rect 403 11 408 18
rect 410 11 415 31
rect 417 25 424 31
rect 452 25 459 31
rect 417 15 426 25
rect 417 13 420 15
rect 422 13 426 15
rect 417 11 426 13
rect 428 22 435 25
rect 428 20 431 22
rect 433 20 435 22
rect 428 18 435 20
rect 441 22 448 25
rect 441 20 443 22
rect 445 20 448 22
rect 441 18 448 20
rect 428 11 433 18
rect 443 11 448 18
rect 450 15 459 25
rect 450 13 454 15
rect 456 13 459 15
rect 450 11 459 13
rect 461 11 466 31
rect 468 24 473 31
rect 479 29 486 31
rect 479 27 481 29
rect 483 27 486 29
rect 468 22 475 24
rect 468 20 471 22
rect 473 20 475 22
rect 468 18 475 20
rect 479 22 486 27
rect 479 20 481 22
rect 483 20 486 22
rect 468 11 473 18
rect 479 17 486 20
rect 488 29 496 31
rect 488 27 491 29
rect 493 27 496 29
rect 488 17 496 27
rect 498 24 503 31
rect 529 24 536 26
rect 498 21 506 24
rect 498 19 501 21
rect 503 19 506 21
rect 498 17 506 19
rect 501 14 506 17
rect 508 18 516 24
rect 508 16 511 18
rect 513 16 516 18
rect 508 14 516 16
rect 511 11 516 14
rect 518 22 525 24
rect 518 20 521 22
rect 523 20 525 22
rect 529 22 531 24
rect 533 22 536 24
rect 529 20 536 22
rect 538 24 546 26
rect 538 22 541 24
rect 543 22 546 24
rect 538 20 546 22
rect 548 24 556 26
rect 548 22 551 24
rect 553 22 556 24
rect 548 20 556 22
rect 558 24 565 26
rect 581 25 588 31
rect 558 22 561 24
rect 563 22 565 24
rect 558 20 565 22
rect 570 22 577 25
rect 570 20 572 22
rect 574 20 577 22
rect 518 18 525 20
rect 518 11 523 18
rect 570 18 577 20
rect 572 11 577 18
rect 579 15 588 25
rect 579 13 583 15
rect 585 13 588 15
rect 579 11 588 13
rect 590 11 595 31
rect 597 24 602 31
rect 608 29 615 31
rect 608 27 610 29
rect 612 27 615 29
rect 597 22 604 24
rect 597 20 600 22
rect 602 20 604 22
rect 597 18 604 20
rect 608 22 615 27
rect 608 20 610 22
rect 612 20 615 22
rect 597 11 602 18
rect 608 17 615 20
rect 617 29 625 31
rect 617 27 620 29
rect 622 27 625 29
rect 617 17 625 27
rect 627 24 632 31
rect 673 25 680 31
rect 627 21 635 24
rect 627 19 630 21
rect 632 19 635 21
rect 627 17 635 19
rect 630 14 635 17
rect 637 18 645 24
rect 637 16 640 18
rect 642 16 645 18
rect 637 14 645 16
rect 640 11 645 14
rect 647 22 654 24
rect 647 20 650 22
rect 652 20 654 22
rect 647 18 654 20
rect 662 22 669 25
rect 662 20 664 22
rect 666 20 669 22
rect 662 18 669 20
rect 647 11 652 18
rect 664 11 669 18
rect 671 15 680 25
rect 671 13 675 15
rect 677 13 680 15
rect 671 11 680 13
rect 682 11 687 31
rect 689 24 694 31
rect 700 29 707 31
rect 700 27 702 29
rect 704 27 707 29
rect 689 22 696 24
rect 689 20 692 22
rect 694 20 696 22
rect 689 18 696 20
rect 700 22 707 27
rect 700 20 702 22
rect 704 20 707 22
rect 689 11 694 18
rect 700 17 707 20
rect 709 29 717 31
rect 709 27 712 29
rect 714 27 717 29
rect 709 17 717 27
rect 719 24 724 31
rect 719 21 727 24
rect 719 19 722 21
rect 724 19 727 21
rect 719 17 727 19
rect 722 14 727 17
rect 729 18 737 24
rect 729 16 732 18
rect 734 16 737 18
rect 729 14 737 16
rect 732 11 737 14
rect 739 22 746 24
rect 739 20 742 22
rect 744 20 746 22
rect 739 18 746 20
rect 739 11 744 18
<< pdif >>
rect 5 56 10 71
rect 3 54 10 56
rect 3 52 5 54
rect 7 52 10 54
rect 3 47 10 52
rect 3 45 5 47
rect 7 45 10 47
rect 3 43 10 45
rect 12 69 20 71
rect 12 67 15 69
rect 17 67 20 69
rect 12 62 20 67
rect 12 60 15 62
rect 17 60 20 62
rect 12 43 20 60
rect 22 61 30 71
rect 22 59 25 61
rect 27 59 30 61
rect 22 54 30 59
rect 22 52 25 54
rect 27 52 30 54
rect 22 43 30 52
rect 32 69 46 71
rect 32 67 37 69
rect 39 68 46 69
rect 69 69 78 71
rect 39 67 48 68
rect 32 62 48 67
rect 32 60 37 62
rect 39 60 48 62
rect 32 43 48 60
rect 50 43 55 68
rect 57 59 62 68
rect 69 67 72 69
rect 74 67 78 69
rect 69 59 78 67
rect 57 50 65 59
rect 57 48 60 50
rect 62 48 65 50
rect 57 46 65 48
rect 67 46 78 59
rect 80 59 85 71
rect 93 64 98 71
rect 91 62 98 64
rect 91 60 93 62
rect 95 60 98 62
rect 80 57 87 59
rect 91 58 98 60
rect 80 55 83 57
rect 85 55 87 57
rect 80 50 87 55
rect 93 53 98 58
rect 100 53 105 71
rect 107 69 116 71
rect 107 67 111 69
rect 113 67 116 69
rect 107 62 116 67
rect 107 53 118 62
rect 80 48 83 50
rect 85 48 87 50
rect 80 46 87 48
rect 57 43 62 46
rect 110 50 118 53
rect 120 60 127 62
rect 120 58 123 60
rect 125 58 127 60
rect 120 56 127 58
rect 134 56 139 71
rect 120 50 125 56
rect 132 54 139 56
rect 132 52 134 54
rect 136 52 139 54
rect 132 47 139 52
rect 132 45 134 47
rect 136 45 139 47
rect 132 43 139 45
rect 141 69 149 71
rect 141 67 144 69
rect 146 67 149 69
rect 141 62 149 67
rect 141 60 144 62
rect 146 60 149 62
rect 141 43 149 60
rect 151 61 159 71
rect 151 59 154 61
rect 156 59 159 61
rect 151 54 159 59
rect 151 52 154 54
rect 156 52 159 54
rect 151 43 159 52
rect 161 69 175 71
rect 161 67 166 69
rect 168 68 175 69
rect 198 69 207 71
rect 168 67 177 68
rect 161 62 177 67
rect 161 60 166 62
rect 168 60 177 62
rect 161 43 177 60
rect 179 43 184 68
rect 186 59 191 68
rect 198 67 201 69
rect 203 67 207 69
rect 198 59 207 67
rect 186 50 194 59
rect 186 48 189 50
rect 191 48 194 50
rect 186 46 194 48
rect 196 46 207 59
rect 209 59 214 71
rect 224 59 229 71
rect 209 57 216 59
rect 209 55 212 57
rect 214 55 216 57
rect 209 50 216 55
rect 209 48 212 50
rect 214 48 216 50
rect 209 46 216 48
rect 222 57 229 59
rect 222 55 224 57
rect 226 55 229 57
rect 222 50 229 55
rect 222 48 224 50
rect 226 48 229 50
rect 222 46 229 48
rect 231 69 240 71
rect 231 67 235 69
rect 237 67 240 69
rect 263 69 277 71
rect 263 68 270 69
rect 231 59 240 67
rect 247 59 252 68
rect 231 46 242 59
rect 244 50 252 59
rect 244 48 247 50
rect 249 48 252 50
rect 244 46 252 48
rect 186 43 191 46
rect 247 43 252 46
rect 254 43 259 68
rect 261 67 270 68
rect 272 67 277 69
rect 261 62 277 67
rect 261 60 270 62
rect 272 60 277 62
rect 261 43 277 60
rect 279 61 287 71
rect 279 59 282 61
rect 284 59 287 61
rect 279 54 287 59
rect 279 52 282 54
rect 284 52 287 54
rect 279 43 287 52
rect 289 69 297 71
rect 289 67 292 69
rect 294 67 297 69
rect 289 62 297 67
rect 289 60 292 62
rect 294 60 297 62
rect 289 43 297 60
rect 299 56 304 71
rect 322 69 331 71
rect 322 67 325 69
rect 327 67 331 69
rect 322 62 331 67
rect 311 60 318 62
rect 311 58 313 60
rect 315 58 318 60
rect 311 56 318 58
rect 299 54 306 56
rect 299 52 302 54
rect 304 52 306 54
rect 299 47 306 52
rect 313 50 318 56
rect 320 53 331 62
rect 333 53 338 71
rect 340 64 345 71
rect 340 62 347 64
rect 340 60 343 62
rect 345 60 347 62
rect 340 58 347 60
rect 353 59 358 71
rect 340 53 345 58
rect 351 57 358 59
rect 351 55 353 57
rect 355 55 358 57
rect 320 50 328 53
rect 299 45 302 47
rect 304 45 306 47
rect 299 43 306 45
rect 351 50 358 55
rect 351 48 353 50
rect 355 48 358 50
rect 351 46 358 48
rect 360 69 369 71
rect 360 67 364 69
rect 366 67 369 69
rect 392 69 406 71
rect 392 68 399 69
rect 360 59 369 67
rect 376 59 381 68
rect 360 46 371 59
rect 373 50 381 59
rect 373 48 376 50
rect 378 48 381 50
rect 373 46 381 48
rect 376 43 381 46
rect 383 43 388 68
rect 390 67 399 68
rect 401 67 406 69
rect 390 62 406 67
rect 390 60 399 62
rect 401 60 406 62
rect 390 43 406 60
rect 408 61 416 71
rect 408 59 411 61
rect 413 59 416 61
rect 408 54 416 59
rect 408 52 411 54
rect 413 52 416 54
rect 408 43 416 52
rect 418 69 426 71
rect 418 67 421 69
rect 423 67 426 69
rect 418 62 426 67
rect 418 60 421 62
rect 423 60 426 62
rect 418 43 426 60
rect 428 56 433 71
rect 443 56 448 71
rect 428 54 435 56
rect 428 52 431 54
rect 433 52 435 54
rect 428 47 435 52
rect 428 45 431 47
rect 433 45 435 47
rect 428 43 435 45
rect 441 54 448 56
rect 441 52 443 54
rect 445 52 448 54
rect 441 47 448 52
rect 441 45 443 47
rect 445 45 448 47
rect 441 43 448 45
rect 450 69 458 71
rect 450 67 453 69
rect 455 67 458 69
rect 450 62 458 67
rect 450 60 453 62
rect 455 60 458 62
rect 450 43 458 60
rect 460 61 468 71
rect 460 59 463 61
rect 465 59 468 61
rect 460 54 468 59
rect 460 52 463 54
rect 465 52 468 54
rect 460 43 468 52
rect 470 69 484 71
rect 470 67 475 69
rect 477 68 484 69
rect 507 69 516 71
rect 477 67 486 68
rect 470 62 486 67
rect 470 60 475 62
rect 477 60 486 62
rect 470 43 486 60
rect 488 43 493 68
rect 495 59 500 68
rect 507 67 510 69
rect 512 67 516 69
rect 507 59 516 67
rect 495 50 503 59
rect 495 48 498 50
rect 500 48 503 50
rect 495 46 503 48
rect 505 46 516 59
rect 518 59 523 71
rect 531 64 536 71
rect 529 62 536 64
rect 529 60 531 62
rect 533 60 536 62
rect 518 57 525 59
rect 529 58 536 60
rect 518 55 521 57
rect 523 55 525 57
rect 518 50 525 55
rect 531 53 536 58
rect 538 53 543 71
rect 545 69 554 71
rect 545 67 549 69
rect 551 67 554 69
rect 545 62 554 67
rect 545 53 556 62
rect 518 48 521 50
rect 523 48 525 50
rect 518 46 525 48
rect 495 43 500 46
rect 548 50 556 53
rect 558 60 565 62
rect 558 58 561 60
rect 563 58 565 60
rect 558 56 565 58
rect 572 56 577 71
rect 558 50 563 56
rect 570 54 577 56
rect 570 52 572 54
rect 574 52 577 54
rect 570 47 577 52
rect 570 45 572 47
rect 574 45 577 47
rect 570 43 577 45
rect 579 69 587 71
rect 579 67 582 69
rect 584 67 587 69
rect 579 62 587 67
rect 579 60 582 62
rect 584 60 587 62
rect 579 43 587 60
rect 589 61 597 71
rect 589 59 592 61
rect 594 59 597 61
rect 589 54 597 59
rect 589 52 592 54
rect 594 52 597 54
rect 589 43 597 52
rect 599 69 613 71
rect 599 67 604 69
rect 606 68 613 69
rect 636 69 645 71
rect 606 67 615 68
rect 599 62 615 67
rect 599 60 604 62
rect 606 60 615 62
rect 599 43 615 60
rect 617 43 622 68
rect 624 59 629 68
rect 636 67 639 69
rect 641 67 645 69
rect 636 59 645 67
rect 624 50 632 59
rect 624 48 627 50
rect 629 48 632 50
rect 624 46 632 48
rect 634 46 645 59
rect 647 59 652 71
rect 647 57 654 59
rect 647 55 650 57
rect 652 55 654 57
rect 664 56 669 71
rect 647 50 654 55
rect 647 48 650 50
rect 652 48 654 50
rect 647 46 654 48
rect 662 54 669 56
rect 662 52 664 54
rect 666 52 669 54
rect 662 47 669 52
rect 624 43 629 46
rect 662 45 664 47
rect 666 45 669 47
rect 662 43 669 45
rect 671 69 679 71
rect 671 67 674 69
rect 676 67 679 69
rect 671 62 679 67
rect 671 60 674 62
rect 676 60 679 62
rect 671 43 679 60
rect 681 61 689 71
rect 681 59 684 61
rect 686 59 689 61
rect 681 54 689 59
rect 681 52 684 54
rect 686 52 689 54
rect 681 43 689 52
rect 691 69 705 71
rect 691 67 696 69
rect 698 68 705 69
rect 728 69 737 71
rect 698 67 707 68
rect 691 62 707 67
rect 691 60 696 62
rect 698 60 707 62
rect 691 43 707 60
rect 709 43 714 68
rect 716 59 721 68
rect 728 67 731 69
rect 733 67 737 69
rect 728 59 737 67
rect 716 50 724 59
rect 716 48 719 50
rect 721 48 724 50
rect 716 46 724 48
rect 726 46 737 59
rect 739 59 744 71
rect 739 57 746 59
rect 739 55 742 57
rect 744 55 746 57
rect 739 50 746 55
rect 739 48 742 50
rect 744 48 746 50
rect 739 46 746 48
rect 716 43 721 46
<< alu1 >>
rect 0 72 751 77
rect 0 70 122 72
rect 124 70 314 72
rect 316 70 560 72
rect 562 70 751 72
rect 0 69 751 70
rect 74 59 87 63
rect 114 60 127 63
rect 114 59 123 60
rect 2 54 8 56
rect 82 57 87 59
rect 82 55 83 57
rect 85 55 87 57
rect 2 52 5 54
rect 7 52 8 54
rect 2 47 8 52
rect 2 45 5 47
rect 7 45 8 47
rect 2 43 8 45
rect 2 23 6 43
rect 18 43 56 47
rect 51 40 56 43
rect 26 38 41 39
rect 26 36 30 38
rect 32 36 37 38
rect 39 36 41 38
rect 26 35 41 36
rect 51 38 59 40
rect 51 36 56 38
rect 58 36 59 38
rect 35 26 39 35
rect 51 34 59 36
rect 82 50 87 55
rect 82 48 83 50
rect 85 48 87 50
rect 82 46 87 48
rect 83 38 87 46
rect 83 36 84 38
rect 86 36 87 38
rect 2 22 24 23
rect 2 20 5 22
rect 7 20 24 22
rect 2 19 24 20
rect 83 24 87 36
rect 91 47 95 48
rect 91 45 92 47
rect 94 45 95 47
rect 91 39 95 45
rect 99 47 103 56
rect 125 58 127 60
rect 203 59 216 63
rect 99 46 112 47
rect 99 44 106 46
rect 108 44 109 46
rect 111 44 112 46
rect 99 43 112 44
rect 91 38 104 39
rect 91 36 96 38
rect 98 36 104 38
rect 91 35 104 36
rect 91 34 95 35
rect 82 22 87 24
rect 82 20 83 22
rect 85 20 87 22
rect 82 18 87 20
rect 123 26 127 58
rect 122 24 127 26
rect 122 22 123 24
rect 125 22 127 24
rect 122 18 127 22
rect 131 54 137 56
rect 211 57 216 59
rect 211 55 212 57
rect 214 55 216 57
rect 131 52 134 54
rect 136 52 137 54
rect 131 47 137 52
rect 131 45 134 47
rect 136 45 137 47
rect 131 43 137 45
rect 131 23 135 43
rect 147 46 185 47
rect 147 44 173 46
rect 175 44 185 46
rect 147 43 185 44
rect 180 40 185 43
rect 155 38 170 39
rect 155 36 159 38
rect 161 36 166 38
rect 168 36 170 38
rect 155 35 170 36
rect 180 38 188 40
rect 180 36 185 38
rect 187 36 188 38
rect 164 29 168 35
rect 180 34 188 36
rect 211 50 216 55
rect 211 48 212 50
rect 214 48 216 50
rect 211 46 216 48
rect 164 27 165 29
rect 167 27 168 29
rect 164 26 168 27
rect 131 22 153 23
rect 131 20 134 22
rect 136 20 153 22
rect 131 19 153 20
rect 212 24 216 46
rect 211 22 216 24
rect 211 20 212 22
rect 214 20 216 22
rect 211 18 216 20
rect 222 59 235 63
rect 311 60 324 63
rect 222 57 227 59
rect 222 55 224 57
rect 226 55 227 57
rect 311 58 313 60
rect 315 59 324 60
rect 351 59 364 63
rect 512 59 525 63
rect 552 60 565 63
rect 552 59 561 60
rect 222 50 227 55
rect 222 48 224 50
rect 226 48 227 50
rect 222 46 227 48
rect 222 24 226 46
rect 253 46 291 47
rect 253 44 271 46
rect 273 44 291 46
rect 253 43 291 44
rect 253 40 258 43
rect 250 38 258 40
rect 250 36 251 38
rect 253 36 258 38
rect 250 34 258 36
rect 268 38 283 39
rect 268 36 270 38
rect 272 36 277 38
rect 279 36 283 38
rect 268 35 283 36
rect 222 22 227 24
rect 270 29 274 35
rect 301 54 307 56
rect 301 52 302 54
rect 304 52 307 54
rect 301 47 307 52
rect 301 45 302 47
rect 304 45 307 47
rect 301 43 307 45
rect 270 27 271 29
rect 273 27 274 29
rect 270 26 274 27
rect 303 23 307 43
rect 222 20 224 22
rect 226 20 227 22
rect 222 18 227 20
rect 285 22 307 23
rect 285 20 302 22
rect 304 20 307 22
rect 285 19 307 20
rect 311 54 315 58
rect 351 57 356 59
rect 311 52 312 54
rect 314 52 315 54
rect 311 26 315 52
rect 335 47 339 56
rect 351 55 353 57
rect 355 55 356 57
rect 351 50 356 55
rect 351 48 353 50
rect 355 48 356 50
rect 326 46 339 47
rect 326 44 327 46
rect 329 44 330 46
rect 332 44 339 46
rect 326 43 339 44
rect 343 47 347 48
rect 343 45 344 47
rect 346 45 347 47
rect 343 39 347 45
rect 334 38 347 39
rect 334 36 340 38
rect 342 36 347 38
rect 334 35 347 36
rect 343 34 347 35
rect 351 46 356 48
rect 351 38 355 46
rect 351 36 352 38
rect 354 36 355 38
rect 382 43 420 47
rect 311 24 316 26
rect 311 22 313 24
rect 315 22 316 24
rect 311 18 316 22
rect 351 24 355 36
rect 382 40 387 43
rect 379 38 387 40
rect 379 36 380 38
rect 382 36 387 38
rect 379 34 387 36
rect 397 38 412 39
rect 397 36 399 38
rect 401 36 406 38
rect 408 36 412 38
rect 397 35 412 36
rect 351 22 356 24
rect 399 26 403 35
rect 430 54 436 56
rect 430 52 431 54
rect 433 52 436 54
rect 430 47 436 52
rect 430 45 431 47
rect 433 45 436 47
rect 430 43 436 45
rect 432 23 436 43
rect 351 20 353 22
rect 355 20 356 22
rect 351 18 356 20
rect 414 22 436 23
rect 414 20 431 22
rect 433 20 436 22
rect 414 19 436 20
rect 440 54 446 56
rect 520 57 525 59
rect 520 55 521 57
rect 523 55 525 57
rect 440 52 443 54
rect 445 52 446 54
rect 440 47 446 52
rect 440 45 443 47
rect 445 45 446 47
rect 440 43 446 45
rect 440 23 444 43
rect 456 43 494 47
rect 489 40 494 43
rect 464 38 479 39
rect 464 36 468 38
rect 470 36 475 38
rect 477 36 479 38
rect 464 35 479 36
rect 489 38 497 40
rect 489 36 494 38
rect 496 36 497 38
rect 473 26 477 35
rect 489 34 497 36
rect 520 50 525 55
rect 520 48 521 50
rect 523 48 525 50
rect 520 46 525 48
rect 521 38 525 46
rect 521 36 522 38
rect 524 36 525 38
rect 440 22 462 23
rect 440 20 443 22
rect 445 20 462 22
rect 440 19 462 20
rect 521 24 525 36
rect 529 47 533 48
rect 529 45 530 47
rect 532 45 533 47
rect 529 39 533 45
rect 537 47 541 56
rect 563 58 565 60
rect 641 59 654 63
rect 733 59 746 63
rect 561 56 565 58
rect 537 46 550 47
rect 537 44 544 46
rect 546 44 547 46
rect 549 44 550 46
rect 537 43 550 44
rect 529 38 542 39
rect 529 36 534 38
rect 536 36 542 38
rect 529 35 542 36
rect 529 34 533 35
rect 561 54 562 56
rect 564 54 565 56
rect 520 22 525 24
rect 520 20 521 22
rect 523 20 525 22
rect 520 18 525 20
rect 561 26 565 54
rect 560 24 565 26
rect 560 22 561 24
rect 563 22 565 24
rect 560 18 565 22
rect 569 54 575 56
rect 649 57 654 59
rect 649 55 650 57
rect 652 55 654 57
rect 569 52 572 54
rect 574 52 575 54
rect 569 47 575 52
rect 569 45 572 47
rect 574 45 575 47
rect 569 43 575 45
rect 569 23 573 43
rect 585 46 623 47
rect 585 44 609 46
rect 611 44 623 46
rect 585 43 623 44
rect 618 40 623 43
rect 593 38 608 39
rect 593 36 597 38
rect 599 36 604 38
rect 606 36 608 38
rect 593 35 608 36
rect 618 38 626 40
rect 618 36 623 38
rect 625 36 626 38
rect 602 29 606 35
rect 618 34 626 36
rect 649 50 654 55
rect 649 48 650 50
rect 652 48 654 50
rect 649 46 654 48
rect 602 27 603 29
rect 605 27 606 29
rect 602 26 606 27
rect 569 22 591 23
rect 569 20 572 22
rect 574 20 591 22
rect 569 19 591 20
rect 650 24 654 46
rect 649 22 654 24
rect 649 20 650 22
rect 652 20 654 22
rect 649 18 654 20
rect 661 54 667 56
rect 741 57 746 59
rect 741 55 742 57
rect 744 55 746 57
rect 661 52 664 54
rect 666 52 667 54
rect 661 47 667 52
rect 661 45 664 47
rect 666 45 667 47
rect 661 43 667 45
rect 661 37 665 43
rect 677 43 715 47
rect 661 35 662 37
rect 664 35 665 37
rect 661 23 665 35
rect 710 40 715 43
rect 685 38 700 39
rect 685 36 689 38
rect 691 36 696 38
rect 698 36 700 38
rect 685 35 700 36
rect 710 38 718 40
rect 710 36 715 38
rect 717 36 718 38
rect 694 26 698 35
rect 710 34 718 36
rect 741 50 746 55
rect 741 48 742 50
rect 744 48 746 50
rect 741 46 746 48
rect 661 22 683 23
rect 661 20 664 22
rect 666 20 683 22
rect 661 19 683 20
rect 742 24 746 46
rect 741 22 746 24
rect 741 20 742 22
rect 744 20 746 22
rect 741 18 746 20
rect 0 12 751 13
rect 0 10 94 12
rect 96 10 122 12
rect 124 10 314 12
rect 316 10 342 12
rect 344 10 532 12
rect 534 10 560 12
rect 562 10 751 12
rect 0 5 751 10
<< alu2 >>
rect 172 59 315 64
rect 4 47 95 48
rect 131 47 137 48
rect 4 45 5 47
rect 7 45 92 47
rect 94 45 95 47
rect 4 44 95 45
rect 108 46 134 47
rect 108 44 109 46
rect 111 45 134 46
rect 136 45 137 47
rect 111 44 137 45
rect 108 43 137 44
rect 172 46 176 59
rect 172 44 173 46
rect 175 44 176 46
rect 172 43 176 44
rect 270 54 274 55
rect 270 52 271 54
rect 273 52 274 54
rect 270 46 274 52
rect 311 54 315 59
rect 549 59 565 61
rect 549 57 550 59
rect 552 57 565 59
rect 549 56 565 57
rect 311 52 312 54
rect 314 52 315 54
rect 561 54 562 56
rect 564 54 565 56
rect 561 52 565 54
rect 608 60 666 66
rect 311 51 315 52
rect 270 44 271 46
rect 273 44 274 46
rect 270 43 274 44
rect 301 47 307 48
rect 343 47 434 48
rect 301 45 302 47
rect 304 46 330 47
rect 304 45 327 46
rect 301 44 327 45
rect 329 44 330 46
rect 343 45 344 47
rect 346 45 431 47
rect 433 45 434 47
rect 343 44 434 45
rect 442 47 533 48
rect 569 47 575 48
rect 442 45 443 47
rect 445 45 530 47
rect 532 45 533 47
rect 442 44 533 45
rect 546 46 572 47
rect 546 44 547 46
rect 549 45 572 46
rect 574 45 575 47
rect 549 44 575 45
rect 301 43 330 44
rect 546 43 575 44
rect 608 46 613 60
rect 608 44 609 46
rect 611 44 613 46
rect 608 43 613 44
rect 82 38 91 39
rect 82 36 84 38
rect 86 36 91 38
rect 82 35 91 36
rect 87 29 91 35
rect 347 38 356 39
rect 347 36 352 38
rect 354 36 356 38
rect 347 35 356 36
rect 520 38 529 39
rect 520 36 522 38
rect 524 36 529 38
rect 520 35 529 36
rect 125 29 168 30
rect 87 27 165 29
rect 167 27 168 29
rect 87 26 168 27
rect 270 29 313 30
rect 347 29 351 35
rect 270 27 271 29
rect 273 27 351 29
rect 270 26 351 27
rect 87 24 129 26
rect 309 24 351 26
rect 525 29 529 35
rect 661 37 665 60
rect 661 35 662 37
rect 664 35 665 37
rect 661 32 665 35
rect 563 29 606 30
rect 525 27 603 29
rect 605 27 606 29
rect 525 26 606 27
rect 525 24 567 26
<< alu3 >>
rect 541 59 553 61
rect 541 57 550 59
rect 552 57 553 59
rect 541 56 553 57
rect 270 54 545 56
rect 270 52 271 54
rect 273 52 545 54
rect 270 51 545 52
<< ptie >>
rect 92 12 126 14
rect 92 10 94 12
rect 96 10 122 12
rect 124 10 126 12
rect 92 8 126 10
rect 312 12 346 14
rect 312 10 314 12
rect 316 10 342 12
rect 344 10 346 12
rect 312 8 346 10
rect 530 12 564 14
rect 530 10 532 12
rect 534 10 560 12
rect 562 10 564 12
rect 530 8 564 10
<< ntie >>
rect 120 72 126 74
rect 120 70 122 72
rect 124 70 126 72
rect 120 68 126 70
rect 312 72 318 74
rect 312 70 314 72
rect 316 70 318 72
rect 312 68 318 70
rect 558 72 564 74
rect 558 70 560 72
rect 562 70 564 72
rect 558 68 564 70
<< nmos >>
rect 10 11 12 25
rect 21 11 23 31
rect 28 11 30 31
rect 48 17 50 31
rect 58 17 60 31
rect 68 14 70 24
rect 78 11 80 24
rect 98 20 100 26
rect 108 20 110 26
rect 118 20 120 26
rect 139 11 141 25
rect 150 11 152 31
rect 157 11 159 31
rect 177 17 179 31
rect 187 17 189 31
rect 197 14 199 24
rect 207 11 209 24
rect 229 11 231 24
rect 239 14 241 24
rect 249 17 251 31
rect 259 17 261 31
rect 279 11 281 31
rect 286 11 288 31
rect 297 11 299 25
rect 318 20 320 26
rect 328 20 330 26
rect 338 20 340 26
rect 358 11 360 24
rect 368 14 370 24
rect 378 17 380 31
rect 388 17 390 31
rect 408 11 410 31
rect 415 11 417 31
rect 426 11 428 25
rect 448 11 450 25
rect 459 11 461 31
rect 466 11 468 31
rect 486 17 488 31
rect 496 17 498 31
rect 506 14 508 24
rect 516 11 518 24
rect 536 20 538 26
rect 546 20 548 26
rect 556 20 558 26
rect 577 11 579 25
rect 588 11 590 31
rect 595 11 597 31
rect 615 17 617 31
rect 625 17 627 31
rect 635 14 637 24
rect 645 11 647 24
rect 669 11 671 25
rect 680 11 682 31
rect 687 11 689 31
rect 707 17 709 31
rect 717 17 719 31
rect 727 14 729 24
rect 737 11 739 24
<< pmos >>
rect 10 43 12 71
rect 20 43 22 71
rect 30 43 32 71
rect 48 43 50 68
rect 55 43 57 68
rect 65 46 67 59
rect 78 46 80 71
rect 98 53 100 71
rect 105 53 107 71
rect 118 50 120 62
rect 139 43 141 71
rect 149 43 151 71
rect 159 43 161 71
rect 177 43 179 68
rect 184 43 186 68
rect 194 46 196 59
rect 207 46 209 71
rect 229 46 231 71
rect 242 46 244 59
rect 252 43 254 68
rect 259 43 261 68
rect 277 43 279 71
rect 287 43 289 71
rect 297 43 299 71
rect 318 50 320 62
rect 331 53 333 71
rect 338 53 340 71
rect 358 46 360 71
rect 371 46 373 59
rect 381 43 383 68
rect 388 43 390 68
rect 406 43 408 71
rect 416 43 418 71
rect 426 43 428 71
rect 448 43 450 71
rect 458 43 460 71
rect 468 43 470 71
rect 486 43 488 68
rect 493 43 495 68
rect 503 46 505 59
rect 516 46 518 71
rect 536 53 538 71
rect 543 53 545 71
rect 556 50 558 62
rect 577 43 579 71
rect 587 43 589 71
rect 597 43 599 71
rect 615 43 617 68
rect 622 43 624 68
rect 632 46 634 59
rect 645 46 647 71
rect 669 43 671 71
rect 679 43 681 71
rect 689 43 691 71
rect 707 43 709 68
rect 714 43 716 68
rect 724 46 726 59
rect 737 46 739 71
<< polyct0 >>
rect 10 36 12 38
rect 20 36 22 38
rect 70 39 72 41
rect 76 29 78 31
rect 116 37 118 39
rect 139 36 141 38
rect 149 36 151 38
rect 199 39 201 41
rect 205 29 207 31
rect 237 39 239 41
rect 231 29 233 31
rect 287 36 289 38
rect 297 36 299 38
rect 320 37 322 39
rect 366 39 368 41
rect 360 29 362 31
rect 416 36 418 38
rect 426 36 428 38
rect 448 36 450 38
rect 458 36 460 38
rect 508 39 510 41
rect 514 29 516 31
rect 554 37 556 39
rect 577 36 579 38
rect 587 36 589 38
rect 637 39 639 41
rect 669 36 671 38
rect 679 36 681 38
rect 643 29 645 31
rect 729 39 731 41
rect 735 29 737 31
<< polyct1 >>
rect 30 36 32 38
rect 37 36 39 38
rect 56 36 58 38
rect 106 44 108 46
rect 96 36 98 38
rect 159 36 161 38
rect 166 36 168 38
rect 185 36 187 38
rect 330 44 332 46
rect 251 36 253 38
rect 270 36 272 38
rect 277 36 279 38
rect 340 36 342 38
rect 380 36 382 38
rect 399 36 401 38
rect 406 36 408 38
rect 468 36 470 38
rect 475 36 477 38
rect 494 36 496 38
rect 544 44 546 46
rect 534 36 536 38
rect 597 36 599 38
rect 604 36 606 38
rect 623 36 625 38
rect 689 36 691 38
rect 696 36 698 38
rect 715 36 717 38
<< ndifct0 >>
rect 16 13 18 15
rect 43 27 45 29
rect 33 20 35 22
rect 43 20 45 22
rect 53 27 55 29
rect 63 19 65 21
rect 73 16 75 18
rect 93 22 95 24
rect 103 22 105 24
rect 113 22 115 24
rect 145 13 147 15
rect 172 27 174 29
rect 162 20 164 22
rect 172 20 174 22
rect 182 27 184 29
rect 192 19 194 21
rect 202 16 204 18
rect 234 16 236 18
rect 244 19 246 21
rect 254 27 256 29
rect 264 27 266 29
rect 264 20 266 22
rect 274 20 276 22
rect 291 13 293 15
rect 323 22 325 24
rect 333 22 335 24
rect 343 22 345 24
rect 363 16 365 18
rect 373 19 375 21
rect 383 27 385 29
rect 393 27 395 29
rect 393 20 395 22
rect 403 20 405 22
rect 420 13 422 15
rect 454 13 456 15
rect 481 27 483 29
rect 471 20 473 22
rect 481 20 483 22
rect 491 27 493 29
rect 501 19 503 21
rect 511 16 513 18
rect 531 22 533 24
rect 541 22 543 24
rect 551 22 553 24
rect 583 13 585 15
rect 610 27 612 29
rect 600 20 602 22
rect 610 20 612 22
rect 620 27 622 29
rect 630 19 632 21
rect 640 16 642 18
rect 675 13 677 15
rect 702 27 704 29
rect 692 20 694 22
rect 702 20 704 22
rect 712 27 714 29
rect 722 19 724 21
rect 732 16 734 18
<< ndifct1 >>
rect 5 20 7 22
rect 83 20 85 22
rect 123 22 125 24
rect 134 20 136 22
rect 212 20 214 22
rect 224 20 226 22
rect 302 20 304 22
rect 313 22 315 24
rect 353 20 355 22
rect 431 20 433 22
rect 443 20 445 22
rect 521 20 523 22
rect 561 22 563 24
rect 572 20 574 22
rect 650 20 652 22
rect 664 20 666 22
rect 742 20 744 22
<< ntiect1 >>
rect 122 70 124 72
rect 314 70 316 72
rect 560 70 562 72
<< ptiect1 >>
rect 94 10 96 12
rect 122 10 124 12
rect 314 10 316 12
rect 342 10 344 12
rect 532 10 534 12
rect 560 10 562 12
<< pdifct0 >>
rect 15 67 17 69
rect 15 60 17 62
rect 25 59 27 61
rect 25 52 27 54
rect 37 67 39 69
rect 37 60 39 62
rect 72 67 74 69
rect 60 48 62 50
rect 93 60 95 62
rect 111 67 113 69
rect 144 67 146 69
rect 144 60 146 62
rect 154 59 156 61
rect 154 52 156 54
rect 166 67 168 69
rect 166 60 168 62
rect 201 67 203 69
rect 189 48 191 50
rect 235 67 237 69
rect 247 48 249 50
rect 270 67 272 69
rect 270 60 272 62
rect 282 59 284 61
rect 282 52 284 54
rect 292 67 294 69
rect 292 60 294 62
rect 325 67 327 69
rect 343 60 345 62
rect 364 67 366 69
rect 376 48 378 50
rect 399 67 401 69
rect 399 60 401 62
rect 411 59 413 61
rect 411 52 413 54
rect 421 67 423 69
rect 421 60 423 62
rect 453 67 455 69
rect 453 60 455 62
rect 463 59 465 61
rect 463 52 465 54
rect 475 67 477 69
rect 475 60 477 62
rect 510 67 512 69
rect 498 48 500 50
rect 531 60 533 62
rect 549 67 551 69
rect 582 67 584 69
rect 582 60 584 62
rect 592 59 594 61
rect 592 52 594 54
rect 604 67 606 69
rect 604 60 606 62
rect 639 67 641 69
rect 627 48 629 50
rect 674 67 676 69
rect 674 60 676 62
rect 684 59 686 61
rect 684 52 686 54
rect 696 67 698 69
rect 696 60 698 62
rect 731 67 733 69
rect 719 48 721 50
<< pdifct1 >>
rect 5 52 7 54
rect 5 45 7 47
rect 83 55 85 57
rect 83 48 85 50
rect 123 58 125 60
rect 134 52 136 54
rect 134 45 136 47
rect 212 55 214 57
rect 212 48 214 50
rect 224 55 226 57
rect 224 48 226 50
rect 313 58 315 60
rect 302 52 304 54
rect 353 55 355 57
rect 302 45 304 47
rect 353 48 355 50
rect 431 52 433 54
rect 431 45 433 47
rect 443 52 445 54
rect 443 45 445 47
rect 521 55 523 57
rect 521 48 523 50
rect 561 58 563 60
rect 572 52 574 54
rect 572 45 574 47
rect 650 55 652 57
rect 650 48 652 50
rect 664 52 666 54
rect 664 45 666 47
rect 742 55 744 57
rect 742 48 744 50
<< alu0 >>
rect 13 67 15 69
rect 17 67 19 69
rect 13 62 19 67
rect 35 67 37 69
rect 39 67 41 69
rect 13 60 15 62
rect 17 60 19 62
rect 13 59 19 60
rect 24 61 28 63
rect 24 59 25 61
rect 27 59 28 61
rect 35 62 41 67
rect 70 67 72 69
rect 74 67 76 69
rect 70 66 76 67
rect 109 67 111 69
rect 113 67 115 69
rect 109 66 115 67
rect 142 67 144 69
rect 146 67 148 69
rect 35 60 37 62
rect 39 60 41 62
rect 35 59 41 60
rect 91 62 111 63
rect 91 60 93 62
rect 95 60 111 62
rect 91 59 111 60
rect 24 55 28 59
rect 47 55 71 59
rect 11 54 51 55
rect 11 52 25 54
rect 27 52 51 54
rect 11 51 51 52
rect 11 40 15 51
rect 59 50 63 52
rect 67 51 73 55
rect 59 48 60 50
rect 62 48 63 50
rect 59 47 63 48
rect 59 43 66 47
rect 9 38 15 40
rect 9 36 10 38
rect 12 36 15 38
rect 9 34 15 36
rect 19 38 23 43
rect 19 36 20 38
rect 22 36 23 38
rect 19 34 23 36
rect 11 31 15 34
rect 11 27 31 31
rect 27 23 31 27
rect 62 32 66 43
rect 69 41 73 51
rect 69 39 70 41
rect 72 39 73 41
rect 69 37 73 39
rect 62 31 80 32
rect 42 29 46 31
rect 62 30 76 31
rect 42 27 43 29
rect 45 27 46 29
rect 27 22 37 23
rect 27 20 33 22
rect 35 20 37 22
rect 27 19 37 20
rect 42 22 46 27
rect 51 29 76 30
rect 78 29 80 31
rect 51 27 53 29
rect 55 28 80 29
rect 55 27 66 28
rect 51 26 66 27
rect 107 55 111 59
rect 122 56 123 59
rect 142 62 148 67
rect 164 67 166 69
rect 168 67 170 69
rect 142 60 144 62
rect 146 60 148 62
rect 142 59 148 60
rect 153 61 157 63
rect 153 59 154 61
rect 156 59 157 61
rect 164 62 170 67
rect 199 67 201 69
rect 203 67 205 69
rect 199 66 205 67
rect 233 67 235 69
rect 237 67 239 69
rect 233 66 239 67
rect 268 67 270 69
rect 272 67 274 69
rect 164 60 166 62
rect 168 60 170 62
rect 164 59 170 60
rect 107 51 119 55
rect 115 39 119 51
rect 115 37 116 39
rect 118 37 119 39
rect 115 32 119 37
rect 102 28 119 32
rect 42 20 43 22
rect 45 21 67 22
rect 45 20 63 21
rect 42 19 63 20
rect 65 19 67 21
rect 42 18 67 19
rect 72 18 76 20
rect 91 24 97 25
rect 91 22 93 24
rect 95 22 97 24
rect 72 16 73 18
rect 75 16 76 18
rect 14 15 20 16
rect 14 13 16 15
rect 18 13 20 15
rect 72 13 76 16
rect 91 13 97 22
rect 102 24 106 28
rect 102 22 103 24
rect 105 22 106 24
rect 102 20 106 22
rect 111 24 117 25
rect 111 22 113 24
rect 115 22 117 24
rect 111 13 117 22
rect 153 55 157 59
rect 176 55 200 59
rect 140 54 180 55
rect 140 52 154 54
rect 156 52 180 54
rect 140 51 180 52
rect 140 40 144 51
rect 188 50 192 52
rect 196 51 202 55
rect 188 48 189 50
rect 191 48 192 50
rect 188 47 192 48
rect 188 43 195 47
rect 138 38 144 40
rect 138 36 139 38
rect 141 36 144 38
rect 138 34 144 36
rect 148 38 152 43
rect 148 36 149 38
rect 151 36 152 38
rect 148 34 152 36
rect 140 31 144 34
rect 140 27 160 31
rect 156 23 160 27
rect 191 32 195 43
rect 198 41 202 51
rect 198 39 199 41
rect 201 39 202 41
rect 198 37 202 39
rect 191 31 209 32
rect 171 29 175 31
rect 191 30 205 31
rect 171 27 172 29
rect 174 27 175 29
rect 156 22 166 23
rect 156 20 162 22
rect 164 20 166 22
rect 156 19 166 20
rect 171 22 175 27
rect 180 29 205 30
rect 207 29 209 31
rect 180 27 182 29
rect 184 28 209 29
rect 184 27 195 28
rect 180 26 195 27
rect 171 20 172 22
rect 174 21 196 22
rect 174 20 192 21
rect 171 19 192 20
rect 194 19 196 21
rect 171 18 196 19
rect 201 18 205 20
rect 268 62 274 67
rect 290 67 292 69
rect 294 67 296 69
rect 268 60 270 62
rect 272 60 274 62
rect 268 59 274 60
rect 281 61 285 63
rect 281 59 282 61
rect 284 59 285 61
rect 290 62 296 67
rect 323 67 325 69
rect 327 67 329 69
rect 323 66 329 67
rect 362 67 364 69
rect 366 67 368 69
rect 362 66 368 67
rect 397 67 399 69
rect 401 67 403 69
rect 290 60 292 62
rect 294 60 296 62
rect 290 59 296 60
rect 238 55 262 59
rect 281 55 285 59
rect 327 62 347 63
rect 327 60 343 62
rect 345 60 347 62
rect 327 59 347 60
rect 397 62 403 67
rect 419 67 421 69
rect 423 67 425 69
rect 397 60 399 62
rect 401 60 403 62
rect 397 59 403 60
rect 410 61 414 63
rect 410 59 411 61
rect 413 59 414 61
rect 419 62 425 67
rect 419 60 421 62
rect 423 60 425 62
rect 419 59 425 60
rect 451 67 453 69
rect 455 67 457 69
rect 451 62 457 67
rect 473 67 475 69
rect 477 67 479 69
rect 451 60 453 62
rect 455 60 457 62
rect 451 59 457 60
rect 462 61 466 63
rect 462 59 463 61
rect 465 59 466 61
rect 473 62 479 67
rect 508 67 510 69
rect 512 67 514 69
rect 508 66 514 67
rect 547 67 549 69
rect 551 67 553 69
rect 547 66 553 67
rect 580 67 582 69
rect 584 67 586 69
rect 473 60 475 62
rect 477 60 479 62
rect 473 59 479 60
rect 529 62 549 63
rect 529 60 531 62
rect 533 60 549 62
rect 529 59 549 60
rect 236 51 242 55
rect 258 54 298 55
rect 258 52 282 54
rect 284 52 298 54
rect 236 41 240 51
rect 246 50 250 52
rect 258 51 298 52
rect 246 48 247 50
rect 249 48 250 50
rect 246 47 250 48
rect 236 39 237 41
rect 239 39 240 41
rect 236 37 240 39
rect 243 43 250 47
rect 243 32 247 43
rect 286 38 290 43
rect 286 36 287 38
rect 289 36 290 38
rect 229 31 247 32
rect 229 29 231 31
rect 233 30 247 31
rect 233 29 258 30
rect 229 28 254 29
rect 243 27 254 28
rect 256 27 258 29
rect 243 26 258 27
rect 263 29 267 31
rect 263 27 264 29
rect 266 27 267 29
rect 263 22 267 27
rect 286 34 290 36
rect 294 40 298 51
rect 294 38 300 40
rect 294 36 297 38
rect 299 36 300 38
rect 294 34 300 36
rect 294 31 298 34
rect 278 27 298 31
rect 278 23 282 27
rect 242 21 264 22
rect 233 18 237 20
rect 242 19 244 21
rect 246 20 264 21
rect 266 20 267 22
rect 246 19 267 20
rect 272 22 282 23
rect 272 20 274 22
rect 276 20 282 22
rect 272 19 282 20
rect 315 56 316 59
rect 327 55 331 59
rect 319 51 331 55
rect 319 39 323 51
rect 367 55 391 59
rect 410 55 414 59
rect 319 37 320 39
rect 322 37 323 39
rect 319 32 323 37
rect 365 51 371 55
rect 387 54 427 55
rect 387 52 411 54
rect 413 52 427 54
rect 365 41 369 51
rect 375 50 379 52
rect 387 51 427 52
rect 375 48 376 50
rect 378 48 379 50
rect 375 47 379 48
rect 365 39 366 41
rect 368 39 369 41
rect 365 37 369 39
rect 372 43 379 47
rect 319 28 336 32
rect 242 18 267 19
rect 321 24 327 25
rect 321 22 323 24
rect 325 22 327 24
rect 201 16 202 18
rect 204 16 205 18
rect 143 15 149 16
rect 143 13 145 15
rect 147 13 149 15
rect 201 13 205 16
rect 233 16 234 18
rect 236 16 237 18
rect 233 13 237 16
rect 289 15 295 16
rect 289 13 291 15
rect 293 13 295 15
rect 321 13 327 22
rect 332 24 336 28
rect 332 22 333 24
rect 335 22 336 24
rect 332 20 336 22
rect 341 24 347 25
rect 341 22 343 24
rect 345 22 347 24
rect 341 13 347 22
rect 372 32 376 43
rect 415 38 419 43
rect 415 36 416 38
rect 418 36 419 38
rect 358 31 376 32
rect 358 29 360 31
rect 362 30 376 31
rect 362 29 387 30
rect 358 28 383 29
rect 372 27 383 28
rect 385 27 387 29
rect 372 26 387 27
rect 392 29 396 31
rect 392 27 393 29
rect 395 27 396 29
rect 392 22 396 27
rect 415 34 419 36
rect 423 40 427 51
rect 423 38 429 40
rect 423 36 426 38
rect 428 36 429 38
rect 423 34 429 36
rect 423 31 427 34
rect 407 27 427 31
rect 407 23 411 27
rect 371 21 393 22
rect 362 18 366 20
rect 371 19 373 21
rect 375 20 393 21
rect 395 20 396 22
rect 375 19 396 20
rect 401 22 411 23
rect 401 20 403 22
rect 405 20 411 22
rect 401 19 411 20
rect 462 55 466 59
rect 485 55 509 59
rect 449 54 489 55
rect 449 52 463 54
rect 465 52 489 54
rect 449 51 489 52
rect 449 40 453 51
rect 497 50 501 52
rect 505 51 511 55
rect 497 48 498 50
rect 500 48 501 50
rect 497 47 501 48
rect 497 43 504 47
rect 447 38 453 40
rect 447 36 448 38
rect 450 36 453 38
rect 447 34 453 36
rect 457 38 461 43
rect 457 36 458 38
rect 460 36 461 38
rect 457 34 461 36
rect 449 31 453 34
rect 449 27 469 31
rect 465 23 469 27
rect 500 32 504 43
rect 507 41 511 51
rect 507 39 508 41
rect 510 39 511 41
rect 507 37 511 39
rect 500 31 518 32
rect 480 29 484 31
rect 500 30 514 31
rect 480 27 481 29
rect 483 27 484 29
rect 465 22 475 23
rect 465 20 471 22
rect 473 20 475 22
rect 465 19 475 20
rect 480 22 484 27
rect 489 29 514 30
rect 516 29 518 31
rect 489 27 491 29
rect 493 28 518 29
rect 493 27 504 28
rect 489 26 504 27
rect 545 55 549 59
rect 560 56 561 59
rect 580 62 586 67
rect 602 67 604 69
rect 606 67 608 69
rect 580 60 582 62
rect 584 60 586 62
rect 580 59 586 60
rect 591 61 595 63
rect 591 59 592 61
rect 594 59 595 61
rect 602 62 608 67
rect 637 67 639 69
rect 641 67 643 69
rect 637 66 643 67
rect 672 67 674 69
rect 676 67 678 69
rect 602 60 604 62
rect 606 60 608 62
rect 602 59 608 60
rect 672 62 678 67
rect 694 67 696 69
rect 698 67 700 69
rect 672 60 674 62
rect 676 60 678 62
rect 672 59 678 60
rect 683 61 687 63
rect 683 59 684 61
rect 686 59 687 61
rect 694 62 700 67
rect 729 67 731 69
rect 733 67 735 69
rect 729 66 735 67
rect 694 60 696 62
rect 698 60 700 62
rect 694 59 700 60
rect 545 51 557 55
rect 553 39 557 51
rect 553 37 554 39
rect 556 37 557 39
rect 553 32 557 37
rect 540 28 557 32
rect 480 20 481 22
rect 483 21 505 22
rect 483 20 501 21
rect 480 19 501 20
rect 503 19 505 21
rect 371 18 396 19
rect 480 18 505 19
rect 510 18 514 20
rect 529 24 535 25
rect 529 22 531 24
rect 533 22 535 24
rect 362 16 363 18
rect 365 16 366 18
rect 510 16 511 18
rect 513 16 514 18
rect 362 13 366 16
rect 418 15 424 16
rect 418 13 420 15
rect 422 13 424 15
rect 452 15 458 16
rect 452 13 454 15
rect 456 13 458 15
rect 510 13 514 16
rect 529 13 535 22
rect 540 24 544 28
rect 540 22 541 24
rect 543 22 544 24
rect 540 20 544 22
rect 549 24 555 25
rect 549 22 551 24
rect 553 22 555 24
rect 549 13 555 22
rect 591 55 595 59
rect 614 55 638 59
rect 578 54 618 55
rect 578 52 592 54
rect 594 52 618 54
rect 578 51 618 52
rect 578 40 582 51
rect 626 50 630 52
rect 634 51 640 55
rect 626 48 627 50
rect 629 48 630 50
rect 626 47 630 48
rect 626 43 633 47
rect 576 38 582 40
rect 576 36 577 38
rect 579 36 582 38
rect 576 34 582 36
rect 586 38 590 43
rect 586 36 587 38
rect 589 36 590 38
rect 586 34 590 36
rect 578 31 582 34
rect 578 27 598 31
rect 594 23 598 27
rect 629 32 633 43
rect 636 41 640 51
rect 636 39 637 41
rect 639 39 640 41
rect 636 37 640 39
rect 629 31 647 32
rect 609 29 613 31
rect 629 30 643 31
rect 609 27 610 29
rect 612 27 613 29
rect 594 22 604 23
rect 594 20 600 22
rect 602 20 604 22
rect 594 19 604 20
rect 609 22 613 27
rect 618 29 643 30
rect 645 29 647 31
rect 618 27 620 29
rect 622 28 647 29
rect 622 27 633 28
rect 618 26 633 27
rect 609 20 610 22
rect 612 21 634 22
rect 612 20 630 21
rect 609 19 630 20
rect 632 19 634 21
rect 609 18 634 19
rect 639 18 643 20
rect 683 55 687 59
rect 706 55 730 59
rect 670 54 710 55
rect 670 52 684 54
rect 686 52 710 54
rect 670 51 710 52
rect 670 40 674 51
rect 718 50 722 52
rect 726 51 732 55
rect 718 48 719 50
rect 721 48 722 50
rect 718 47 722 48
rect 718 43 725 47
rect 668 38 674 40
rect 668 36 669 38
rect 671 36 674 38
rect 668 34 674 36
rect 678 38 682 43
rect 678 36 679 38
rect 681 36 682 38
rect 678 34 682 36
rect 670 31 674 34
rect 670 27 690 31
rect 686 23 690 27
rect 721 32 725 43
rect 728 41 732 51
rect 728 39 729 41
rect 731 39 732 41
rect 728 37 732 39
rect 721 31 739 32
rect 701 29 705 31
rect 721 30 735 31
rect 701 27 702 29
rect 704 27 705 29
rect 686 22 696 23
rect 686 20 692 22
rect 694 20 696 22
rect 686 19 696 20
rect 701 22 705 27
rect 710 29 735 30
rect 737 29 739 31
rect 710 27 712 29
rect 714 28 739 29
rect 714 27 725 28
rect 710 26 725 27
rect 701 20 702 22
rect 704 21 726 22
rect 704 20 722 21
rect 701 19 722 20
rect 724 19 726 21
rect 701 18 726 19
rect 731 18 735 20
rect 639 16 640 18
rect 642 16 643 18
rect 731 16 732 18
rect 734 16 735 18
rect 581 15 587 16
rect 581 13 583 15
rect 585 13 587 15
rect 639 13 643 16
rect 673 15 679 16
rect 673 13 675 15
rect 677 13 679 15
rect 731 13 735 16
<< via1 >>
rect 5 45 7 47
rect 84 36 86 38
rect 92 45 94 47
rect 109 44 111 46
rect 134 45 136 47
rect 173 44 175 46
rect 165 27 167 29
rect 271 44 273 46
rect 302 45 304 47
rect 271 27 273 29
rect 312 52 314 54
rect 327 44 329 46
rect 344 45 346 47
rect 352 36 354 38
rect 431 45 433 47
rect 443 45 445 47
rect 522 36 524 38
rect 530 45 532 47
rect 547 44 549 46
rect 562 54 564 56
rect 572 45 574 47
rect 609 44 611 46
rect 603 27 605 29
rect 662 35 664 37
<< via2 >>
rect 271 52 273 54
rect 550 57 552 59
<< labels >>
rlabel alu1 170 73 170 73 4 vdd
rlabel alu1 170 9 170 9 4 vss
rlabel alu1 37 33 37 33 1 a4
rlabel alu1 53 38 53 38 1 b4
rlabel alu1 158 45 158 45 1 ci4
rlabel alu1 214 37 214 37 1 so4
rlabel alu1 224 37 224 37 1 so3
rlabel alu1 280 45 280 45 1 ci3
rlabel alu1 125 37 125 37 1 co4
rlabel alu1 313 37 313 37 1 co3
rlabel alu1 563 37 563 37 1 co2
rlabel alu1 652 37 652 37 1 so2
rlabel alu1 596 45 596 45 1 ci2
rlabel alu1 475 33 475 33 1 a2
rlabel alu1 401 33 401 33 1 a3
rlabel alu1 385 37 385 37 1 b3
rlabel alu1 491 37 491 37 1 b2
rlabel alu1 744 37 744 37 1 so1
rlabel alu2 664 49 664 49 1 co1
rlabel alu1 688 37 688 37 1 a1
rlabel alu1 680 45 680 45 1 b1
<< end >>
