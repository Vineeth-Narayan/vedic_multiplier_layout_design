magic
tech scmos
timestamp 1636138048
<< ab >>
rect 6 101 46 173
rect 49 160 89 173
rect 49 156 74 160
rect 58 154 74 156
rect 79 154 89 160
rect 58 152 89 154
rect 49 101 89 152
rect 92 160 132 173
rect 92 152 109 160
rect 122 154 132 160
rect 117 152 132 154
rect 92 101 132 152
rect 135 101 175 173
rect 5 5 97 77
rect 99 5 197 77
<< nwell >>
rect 4 133 177 178
rect 3 37 197 82
<< pwell >>
rect 4 96 177 133
rect 3 0 197 37
<< poly >>
rect 46 160 72 162
rect 78 160 158 162
rect 25 158 31 160
rect 25 156 27 158
rect 29 156 31 158
rect 15 151 17 156
rect 25 154 31 156
rect 46 154 48 160
rect 68 158 74 160
rect 68 156 70 158
rect 72 156 74 158
rect 25 149 27 154
rect 35 152 48 154
rect 35 149 37 152
rect 58 151 60 156
rect 68 154 74 156
rect 68 149 70 154
rect 78 149 80 160
rect 154 158 160 160
rect 154 156 156 158
rect 158 156 160 158
rect 101 151 103 156
rect 111 149 113 153
rect 121 149 123 154
rect 144 151 146 156
rect 154 154 160 156
rect 154 149 156 154
rect 164 149 166 154
rect 15 136 17 139
rect 25 136 27 139
rect 15 134 21 136
rect 15 132 17 134
rect 19 132 21 134
rect 25 133 29 136
rect 15 130 21 132
rect 15 122 17 130
rect 27 119 29 133
rect 35 128 37 139
rect 58 136 60 139
rect 68 136 70 139
rect 58 134 64 136
rect 58 132 60 134
rect 62 132 64 134
rect 68 133 72 136
rect 58 130 64 132
rect 34 126 40 128
rect 34 124 36 126
rect 38 124 40 126
rect 34 122 40 124
rect 58 122 60 130
rect 34 119 36 122
rect 15 112 17 116
rect 70 119 72 133
rect 78 128 80 139
rect 101 136 103 139
rect 111 136 113 139
rect 101 134 107 136
rect 101 132 103 134
rect 105 132 107 134
rect 111 133 115 136
rect 101 130 107 132
rect 77 126 83 128
rect 77 124 79 126
rect 81 124 83 126
rect 77 122 83 124
rect 101 122 103 130
rect 77 119 79 122
rect 58 112 60 116
rect 113 119 115 133
rect 121 128 123 139
rect 144 136 146 139
rect 154 136 156 139
rect 144 134 150 136
rect 144 132 146 134
rect 148 132 150 134
rect 154 133 158 136
rect 144 130 150 132
rect 120 126 126 128
rect 120 124 122 126
rect 124 124 126 126
rect 120 122 126 124
rect 144 122 146 130
rect 120 119 122 122
rect 101 112 103 116
rect 156 119 158 133
rect 164 128 166 139
rect 163 126 169 128
rect 163 124 165 126
rect 167 124 169 126
rect 163 122 169 124
rect 163 119 165 122
rect 144 112 146 116
rect 27 98 29 110
rect 34 105 36 110
rect 70 105 72 110
rect 77 105 79 110
rect 113 98 115 110
rect 120 98 122 110
rect 156 105 158 110
rect 163 98 165 110
rect 27 96 116 98
rect 120 96 165 98
rect 14 71 16 75
rect 37 68 39 73
rect 44 68 46 73
rect 62 71 64 75
rect 72 71 74 75
rect 82 71 84 75
rect 116 71 118 75
rect 126 71 128 75
rect 136 71 138 75
rect 27 59 29 64
rect 14 33 16 46
rect 27 43 29 46
rect 154 68 156 73
rect 161 68 163 73
rect 184 71 186 75
rect 171 59 173 64
rect 171 43 173 46
rect 20 41 29 43
rect 20 39 22 41
rect 24 39 26 41
rect 37 40 39 43
rect 44 40 46 43
rect 62 40 64 43
rect 72 40 74 43
rect 82 40 84 43
rect 116 40 118 43
rect 126 40 128 43
rect 136 40 138 43
rect 154 40 156 43
rect 161 40 163 43
rect 171 41 180 43
rect 20 37 26 39
rect 14 31 20 33
rect 14 29 16 31
rect 18 29 20 31
rect 14 27 20 29
rect 14 24 16 27
rect 24 24 26 37
rect 34 38 40 40
rect 34 36 36 38
rect 38 36 40 38
rect 34 34 40 36
rect 44 38 66 40
rect 44 36 55 38
rect 57 36 62 38
rect 64 36 66 38
rect 44 34 66 36
rect 70 38 76 40
rect 70 36 72 38
rect 74 36 76 38
rect 70 34 76 36
rect 80 38 86 40
rect 80 36 82 38
rect 84 36 86 38
rect 80 34 86 36
rect 114 38 120 40
rect 114 36 116 38
rect 118 36 120 38
rect 114 34 120 36
rect 124 38 130 40
rect 124 36 126 38
rect 128 36 130 38
rect 124 34 130 36
rect 134 38 156 40
rect 134 36 136 38
rect 138 36 143 38
rect 145 36 156 38
rect 134 34 156 36
rect 160 38 166 40
rect 160 36 162 38
rect 164 36 166 38
rect 160 34 166 36
rect 34 31 36 34
rect 44 31 46 34
rect 64 31 66 34
rect 71 31 73 34
rect 14 7 16 11
rect 24 9 26 14
rect 34 12 36 17
rect 44 12 46 17
rect 82 25 84 34
rect 116 25 118 34
rect 127 31 129 34
rect 134 31 136 34
rect 154 31 156 34
rect 164 31 166 34
rect 174 39 176 41
rect 178 39 180 41
rect 174 37 180 39
rect 174 24 176 37
rect 184 33 186 46
rect 180 31 186 33
rect 180 29 182 31
rect 184 29 186 31
rect 180 27 186 29
rect 184 24 186 27
rect 154 12 156 17
rect 164 12 166 17
rect 64 7 66 11
rect 71 7 73 11
rect 82 7 84 11
rect 116 7 118 11
rect 127 7 129 11
rect 134 7 136 11
rect 174 9 176 14
rect 184 7 186 11
<< ndif >>
rect 8 120 15 122
rect 8 118 10 120
rect 12 118 15 120
rect 8 116 15 118
rect 17 119 25 122
rect 51 120 58 122
rect 17 116 27 119
rect 19 110 27 116
rect 29 110 34 119
rect 36 117 43 119
rect 36 115 39 117
rect 41 115 43 117
rect 51 118 53 120
rect 55 118 58 120
rect 51 116 58 118
rect 60 119 68 122
rect 94 120 101 122
rect 60 116 70 119
rect 36 113 43 115
rect 36 110 41 113
rect 62 110 70 116
rect 72 110 77 119
rect 79 117 86 119
rect 79 115 82 117
rect 84 115 86 117
rect 94 118 96 120
rect 98 118 101 120
rect 94 116 101 118
rect 103 119 111 122
rect 137 120 144 122
rect 103 116 113 119
rect 79 113 86 115
rect 79 110 84 113
rect 105 110 113 116
rect 115 110 120 119
rect 122 117 129 119
rect 122 115 125 117
rect 127 115 129 117
rect 137 118 139 120
rect 141 118 144 120
rect 137 116 144 118
rect 146 119 154 122
rect 146 116 156 119
rect 122 113 129 115
rect 122 110 127 113
rect 148 110 156 116
rect 158 110 163 119
rect 165 117 172 119
rect 165 115 168 117
rect 170 115 172 117
rect 165 113 172 115
rect 165 110 170 113
rect 19 108 25 110
rect 19 106 21 108
rect 23 106 25 108
rect 19 104 25 106
rect 62 108 68 110
rect 62 106 64 108
rect 66 106 68 108
rect 62 104 68 106
rect 105 108 111 110
rect 105 106 107 108
rect 109 106 111 108
rect 105 104 111 106
rect 148 108 154 110
rect 148 106 150 108
rect 152 106 154 108
rect 148 104 154 106
rect 29 24 34 31
rect 7 22 14 24
rect 7 20 9 22
rect 11 20 14 22
rect 7 18 14 20
rect 9 11 14 18
rect 16 18 24 24
rect 16 16 19 18
rect 21 16 24 18
rect 16 14 24 16
rect 26 21 34 24
rect 26 19 29 21
rect 31 19 34 21
rect 26 17 34 19
rect 36 29 44 31
rect 36 27 39 29
rect 41 27 44 29
rect 36 17 44 27
rect 46 29 53 31
rect 46 27 49 29
rect 51 27 53 29
rect 46 22 53 27
rect 59 24 64 31
rect 46 20 49 22
rect 51 20 53 22
rect 46 17 53 20
rect 57 22 64 24
rect 57 20 59 22
rect 61 20 64 22
rect 57 18 64 20
rect 26 14 31 17
rect 16 11 21 14
rect 59 11 64 18
rect 66 11 71 31
rect 73 25 80 31
rect 120 25 127 31
rect 73 15 82 25
rect 73 13 76 15
rect 78 13 82 15
rect 73 11 82 13
rect 84 22 91 25
rect 84 20 87 22
rect 89 20 91 22
rect 84 18 91 20
rect 109 22 116 25
rect 109 20 111 22
rect 113 20 116 22
rect 109 18 116 20
rect 84 11 89 18
rect 111 11 116 18
rect 118 15 127 25
rect 118 13 122 15
rect 124 13 127 15
rect 118 11 127 13
rect 129 11 134 31
rect 136 24 141 31
rect 147 29 154 31
rect 147 27 149 29
rect 151 27 154 29
rect 136 22 143 24
rect 136 20 139 22
rect 141 20 143 22
rect 136 18 143 20
rect 147 22 154 27
rect 147 20 149 22
rect 151 20 154 22
rect 136 11 141 18
rect 147 17 154 20
rect 156 29 164 31
rect 156 27 159 29
rect 161 27 164 29
rect 156 17 164 27
rect 166 24 171 31
rect 166 21 174 24
rect 166 19 169 21
rect 171 19 174 21
rect 166 17 174 19
rect 169 14 174 17
rect 176 18 184 24
rect 176 16 179 18
rect 181 16 184 18
rect 176 14 184 16
rect 179 11 184 14
rect 186 22 193 24
rect 186 20 189 22
rect 191 20 193 22
rect 186 18 193 20
rect 186 11 191 18
<< pdif >>
rect 10 145 15 151
rect 8 143 15 145
rect 8 141 10 143
rect 12 141 15 143
rect 8 139 15 141
rect 17 149 23 151
rect 17 143 25 149
rect 17 141 20 143
rect 22 141 25 143
rect 17 139 25 141
rect 27 143 35 149
rect 27 141 30 143
rect 32 141 35 143
rect 27 139 35 141
rect 37 147 44 149
rect 37 145 40 147
rect 42 145 44 147
rect 53 145 58 151
rect 37 139 44 145
rect 51 143 58 145
rect 51 141 53 143
rect 55 141 58 143
rect 51 139 58 141
rect 60 149 66 151
rect 60 143 68 149
rect 60 141 63 143
rect 65 141 68 143
rect 60 139 68 141
rect 70 143 78 149
rect 70 141 73 143
rect 75 141 78 143
rect 70 139 78 141
rect 80 147 87 149
rect 80 145 83 147
rect 85 145 87 147
rect 96 145 101 151
rect 80 139 87 145
rect 94 143 101 145
rect 94 141 96 143
rect 98 141 101 143
rect 94 139 101 141
rect 103 149 109 151
rect 103 143 111 149
rect 103 141 106 143
rect 108 141 111 143
rect 103 139 111 141
rect 113 143 121 149
rect 113 141 116 143
rect 118 141 121 143
rect 113 139 121 141
rect 123 147 130 149
rect 123 145 126 147
rect 128 145 130 147
rect 139 145 144 151
rect 123 139 130 145
rect 137 143 144 145
rect 137 141 139 143
rect 141 141 144 143
rect 137 139 144 141
rect 146 149 152 151
rect 146 143 154 149
rect 146 141 149 143
rect 151 141 154 143
rect 146 139 154 141
rect 156 143 164 149
rect 156 141 159 143
rect 161 141 164 143
rect 156 139 164 141
rect 166 147 173 149
rect 166 145 169 147
rect 171 145 173 147
rect 166 139 173 145
rect 9 59 14 71
rect 7 57 14 59
rect 7 55 9 57
rect 11 55 14 57
rect 7 50 14 55
rect 7 48 9 50
rect 11 48 14 50
rect 7 46 14 48
rect 16 69 25 71
rect 16 67 20 69
rect 22 67 25 69
rect 48 69 62 71
rect 48 68 55 69
rect 16 59 25 67
rect 32 59 37 68
rect 16 46 27 59
rect 29 50 37 59
rect 29 48 32 50
rect 34 48 37 50
rect 29 46 37 48
rect 32 43 37 46
rect 39 43 44 68
rect 46 67 55 68
rect 57 67 62 69
rect 46 62 62 67
rect 46 60 55 62
rect 57 60 62 62
rect 46 43 62 60
rect 64 61 72 71
rect 64 59 67 61
rect 69 59 72 61
rect 64 54 72 59
rect 64 52 67 54
rect 69 52 72 54
rect 64 43 72 52
rect 74 69 82 71
rect 74 67 77 69
rect 79 67 82 69
rect 74 62 82 67
rect 74 60 77 62
rect 79 60 82 62
rect 74 43 82 60
rect 84 56 89 71
rect 111 56 116 71
rect 84 54 91 56
rect 84 52 87 54
rect 89 52 91 54
rect 84 47 91 52
rect 84 45 87 47
rect 89 45 91 47
rect 84 43 91 45
rect 109 54 116 56
rect 109 52 111 54
rect 113 52 116 54
rect 109 47 116 52
rect 109 45 111 47
rect 113 45 116 47
rect 109 43 116 45
rect 118 69 126 71
rect 118 67 121 69
rect 123 67 126 69
rect 118 62 126 67
rect 118 60 121 62
rect 123 60 126 62
rect 118 43 126 60
rect 128 61 136 71
rect 128 59 131 61
rect 133 59 136 61
rect 128 54 136 59
rect 128 52 131 54
rect 133 52 136 54
rect 128 43 136 52
rect 138 69 152 71
rect 138 67 143 69
rect 145 68 152 69
rect 175 69 184 71
rect 145 67 154 68
rect 138 62 154 67
rect 138 60 143 62
rect 145 60 154 62
rect 138 43 154 60
rect 156 43 161 68
rect 163 59 168 68
rect 175 67 178 69
rect 180 67 184 69
rect 175 59 184 67
rect 163 50 171 59
rect 163 48 166 50
rect 168 48 171 50
rect 163 46 171 48
rect 173 46 184 59
rect 186 59 191 71
rect 186 57 193 59
rect 186 55 189 57
rect 191 55 193 57
rect 186 50 193 55
rect 186 48 189 50
rect 191 48 193 50
rect 186 46 193 48
rect 163 43 168 46
<< alu1 >>
rect 4 168 177 173
rect 4 166 11 168
rect 13 166 25 168
rect 27 166 39 168
rect 41 166 54 168
rect 56 166 68 168
rect 70 166 82 168
rect 84 166 97 168
rect 99 166 111 168
rect 113 166 125 168
rect 127 166 140 168
rect 142 166 154 168
rect 156 166 168 168
rect 170 166 177 168
rect 4 165 177 166
rect 8 143 12 152
rect 8 141 10 143
rect 8 127 12 141
rect 23 158 36 160
rect 23 156 27 158
rect 29 156 36 158
rect 23 154 36 156
rect 23 147 29 154
rect 51 143 55 152
rect 51 141 53 143
rect 8 125 9 127
rect 11 125 12 127
rect 8 120 12 125
rect 8 118 10 120
rect 12 118 20 120
rect 8 114 20 118
rect 40 127 44 136
rect 31 126 44 127
rect 31 124 36 126
rect 38 124 44 126
rect 31 122 44 124
rect 51 126 55 141
rect 66 158 74 160
rect 66 156 70 158
rect 72 156 74 158
rect 66 154 74 156
rect 66 147 72 154
rect 94 143 98 152
rect 94 141 96 143
rect 51 124 52 126
rect 54 124 55 126
rect 51 120 55 124
rect 51 118 53 120
rect 55 118 63 120
rect 51 114 63 118
rect 83 127 87 136
rect 74 126 87 127
rect 74 124 79 126
rect 81 124 87 126
rect 74 122 87 124
rect 94 126 98 141
rect 109 147 115 152
rect 137 143 141 152
rect 137 141 139 143
rect 94 124 95 126
rect 97 124 98 126
rect 94 120 98 124
rect 94 118 96 120
rect 98 118 106 120
rect 94 114 106 118
rect 126 127 130 136
rect 117 126 130 127
rect 117 124 122 126
rect 124 124 130 126
rect 117 122 130 124
rect 137 120 141 141
rect 152 158 165 160
rect 152 156 156 158
rect 158 156 165 158
rect 152 154 165 156
rect 152 147 158 154
rect 137 118 139 120
rect 141 118 149 120
rect 137 114 149 118
rect 169 127 173 136
rect 160 126 173 127
rect 160 124 165 126
rect 167 124 173 126
rect 160 122 173 124
rect 4 108 177 109
rect 4 106 11 108
rect 13 106 21 108
rect 23 106 54 108
rect 56 106 64 108
rect 66 106 97 108
rect 99 106 107 108
rect 109 106 140 108
rect 142 106 150 108
rect 152 106 177 108
rect 4 101 177 106
rect 3 69 197 77
rect 7 59 20 63
rect 180 59 193 63
rect 7 57 12 59
rect 7 55 9 57
rect 11 55 12 57
rect 7 50 12 55
rect 7 48 9 50
rect 11 48 12 50
rect 7 46 12 48
rect 7 24 11 46
rect 38 46 76 47
rect 38 44 48 46
rect 50 44 76 46
rect 38 43 76 44
rect 38 40 43 43
rect 35 38 43 40
rect 35 36 36 38
rect 38 36 43 38
rect 35 34 43 36
rect 53 38 68 39
rect 53 36 55 38
rect 57 36 62 38
rect 64 36 68 38
rect 53 35 68 36
rect 55 34 59 35
rect 86 54 92 56
rect 86 52 87 54
rect 89 52 92 54
rect 86 47 92 52
rect 86 45 87 47
rect 89 45 92 47
rect 86 43 92 45
rect 55 32 56 34
rect 58 32 59 34
rect 7 22 12 24
rect 55 26 59 32
rect 88 23 92 43
rect 7 20 9 22
rect 11 20 12 22
rect 7 18 12 20
rect 70 22 92 23
rect 70 20 87 22
rect 89 20 92 22
rect 70 19 92 20
rect 108 54 114 56
rect 188 57 193 59
rect 188 55 189 57
rect 191 55 193 57
rect 108 52 111 54
rect 113 52 114 54
rect 108 47 114 52
rect 108 45 111 47
rect 113 45 114 47
rect 108 43 114 45
rect 108 35 112 43
rect 124 46 162 47
rect 124 44 158 46
rect 160 44 162 46
rect 124 43 162 44
rect 108 33 109 35
rect 111 33 112 35
rect 157 40 162 43
rect 132 38 147 39
rect 132 36 136 38
rect 138 36 143 38
rect 145 36 147 38
rect 132 35 147 36
rect 157 38 165 40
rect 157 36 162 38
rect 164 36 165 38
rect 108 23 112 33
rect 141 26 145 35
rect 157 34 165 36
rect 188 50 193 55
rect 188 48 189 50
rect 191 48 193 50
rect 188 46 193 48
rect 108 22 130 23
rect 108 20 111 22
rect 113 20 130 22
rect 108 19 130 20
rect 189 24 193 46
rect 188 22 193 24
rect 188 20 189 22
rect 191 20 193 22
rect 188 18 193 20
rect 3 5 197 13
<< alu2 >>
rect -1 127 12 128
rect -1 125 9 127
rect 11 125 12 127
rect -1 124 12 125
rect 45 126 55 127
rect 45 124 52 126
rect 54 124 55 126
rect -1 88 4 124
rect 45 123 55 124
rect 88 126 98 127
rect 88 124 95 126
rect 97 124 98 126
rect 88 123 98 124
rect 45 97 50 123
rect 45 92 81 97
rect -1 83 52 88
rect 47 46 52 83
rect 74 85 81 92
rect 88 95 93 123
rect 88 91 162 95
rect 74 79 142 85
rect 47 44 48 46
rect 50 44 52 46
rect 47 43 52 44
rect 134 38 140 79
rect 156 46 162 91
rect 156 44 158 46
rect 160 44 162 46
rect 156 43 162 44
rect 134 36 136 38
rect 138 36 140 38
rect 55 35 112 36
rect 55 34 109 35
rect 55 32 56 34
rect 58 33 109 34
rect 111 33 112 35
rect 134 34 140 36
rect 58 32 112 33
rect 55 31 112 32
<< ptie >>
rect 9 108 15 110
rect 9 106 11 108
rect 13 106 15 108
rect 9 104 15 106
rect 52 108 58 110
rect 52 106 54 108
rect 56 106 58 108
rect 52 104 58 106
rect 95 108 101 110
rect 95 106 97 108
rect 99 106 101 108
rect 95 104 101 106
rect 138 108 144 110
rect 138 106 140 108
rect 142 106 144 108
rect 138 104 144 106
<< ntie >>
rect 9 168 43 170
rect 9 166 11 168
rect 13 166 25 168
rect 27 166 39 168
rect 41 166 43 168
rect 9 164 43 166
rect 52 168 86 170
rect 52 166 54 168
rect 56 166 68 168
rect 70 166 82 168
rect 84 166 86 168
rect 52 164 86 166
rect 95 168 129 170
rect 95 166 97 168
rect 99 166 111 168
rect 113 166 125 168
rect 127 166 129 168
rect 95 164 129 166
rect 138 168 172 170
rect 138 166 140 168
rect 142 166 154 168
rect 156 166 168 168
rect 170 166 172 168
rect 138 164 172 166
<< nmos >>
rect 15 116 17 122
rect 27 110 29 119
rect 34 110 36 119
rect 58 116 60 122
rect 70 110 72 119
rect 77 110 79 119
rect 101 116 103 122
rect 113 110 115 119
rect 120 110 122 119
rect 144 116 146 122
rect 156 110 158 119
rect 163 110 165 119
rect 14 11 16 24
rect 24 14 26 24
rect 34 17 36 31
rect 44 17 46 31
rect 64 11 66 31
rect 71 11 73 31
rect 82 11 84 25
rect 116 11 118 25
rect 127 11 129 31
rect 134 11 136 31
rect 154 17 156 31
rect 164 17 166 31
rect 174 14 176 24
rect 184 11 186 24
<< pmos >>
rect 15 139 17 151
rect 25 139 27 149
rect 35 139 37 149
rect 58 139 60 151
rect 68 139 70 149
rect 78 139 80 149
rect 101 139 103 151
rect 111 139 113 149
rect 121 139 123 149
rect 144 139 146 151
rect 154 139 156 149
rect 164 139 166 149
rect 14 46 16 71
rect 27 46 29 59
rect 37 43 39 68
rect 44 43 46 68
rect 62 43 64 71
rect 72 43 74 71
rect 82 43 84 71
rect 116 43 118 71
rect 126 43 128 71
rect 136 43 138 71
rect 154 43 156 68
rect 161 43 163 68
rect 171 46 173 59
rect 184 46 186 71
<< polyct0 >>
rect 17 132 19 134
rect 60 132 62 134
rect 103 132 105 134
rect 146 132 148 134
rect 22 39 24 41
rect 16 29 18 31
rect 72 36 74 38
rect 82 36 84 38
rect 116 36 118 38
rect 126 36 128 38
rect 176 39 178 41
rect 182 29 184 31
<< polyct1 >>
rect 27 156 29 158
rect 70 156 72 158
rect 156 156 158 158
rect 36 124 38 126
rect 79 124 81 126
rect 122 124 124 126
rect 165 124 167 126
rect 36 36 38 38
rect 55 36 57 38
rect 62 36 64 38
rect 136 36 138 38
rect 143 36 145 38
rect 162 36 164 38
<< ndifct0 >>
rect 39 115 41 117
rect 82 115 84 117
rect 125 115 127 117
rect 168 115 170 117
rect 19 16 21 18
rect 29 19 31 21
rect 39 27 41 29
rect 49 27 51 29
rect 49 20 51 22
rect 59 20 61 22
rect 76 13 78 15
rect 122 13 124 15
rect 149 27 151 29
rect 139 20 141 22
rect 149 20 151 22
rect 159 27 161 29
rect 169 19 171 21
rect 179 16 181 18
<< ndifct1 >>
rect 10 118 12 120
rect 53 118 55 120
rect 96 118 98 120
rect 139 118 141 120
rect 21 106 23 108
rect 64 106 66 108
rect 107 106 109 108
rect 150 106 152 108
rect 9 20 11 22
rect 87 20 89 22
rect 111 20 113 22
rect 189 20 191 22
<< ntiect1 >>
rect 11 166 13 168
rect 25 166 27 168
rect 39 166 41 168
rect 54 166 56 168
rect 68 166 70 168
rect 82 166 84 168
rect 97 166 99 168
rect 111 166 113 168
rect 125 166 127 168
rect 140 166 142 168
rect 154 166 156 168
rect 168 166 170 168
<< ptiect1 >>
rect 11 106 13 108
rect 54 106 56 108
rect 97 106 99 108
rect 140 106 142 108
<< pdifct0 >>
rect 20 141 22 143
rect 30 141 32 143
rect 40 145 42 147
rect 63 141 65 143
rect 73 141 75 143
rect 83 145 85 147
rect 106 141 108 143
rect 116 141 118 143
rect 126 145 128 147
rect 149 141 151 143
rect 159 141 161 143
rect 169 145 171 147
rect 20 67 22 69
rect 32 48 34 50
rect 55 67 57 69
rect 55 60 57 62
rect 67 59 69 61
rect 67 52 69 54
rect 77 67 79 69
rect 77 60 79 62
rect 121 67 123 69
rect 121 60 123 62
rect 131 59 133 61
rect 131 52 133 54
rect 143 67 145 69
rect 143 60 145 62
rect 178 67 180 69
rect 166 48 168 50
<< pdifct1 >>
rect 10 141 12 143
rect 53 141 55 143
rect 96 141 98 143
rect 139 141 141 143
rect 9 55 11 57
rect 9 48 11 50
rect 87 52 89 54
rect 87 45 89 47
rect 111 52 113 54
rect 111 45 113 47
rect 189 55 191 57
rect 189 48 191 50
<< alu0 >>
rect 12 139 13 145
rect 16 144 20 165
rect 39 147 43 165
rect 39 145 40 147
rect 42 145 43 147
rect 16 143 24 144
rect 16 141 20 143
rect 22 141 24 143
rect 16 140 24 141
rect 28 143 34 144
rect 39 143 43 145
rect 28 141 30 143
rect 32 141 34 143
rect 28 135 34 141
rect 15 134 34 135
rect 15 132 17 134
rect 19 132 34 134
rect 15 131 34 132
rect 12 120 13 122
rect 24 118 28 131
rect 55 139 56 145
rect 59 144 63 165
rect 82 147 86 165
rect 82 145 83 147
rect 85 145 86 147
rect 59 143 67 144
rect 59 141 63 143
rect 65 141 67 143
rect 59 140 67 141
rect 71 143 77 144
rect 82 143 86 145
rect 71 141 73 143
rect 75 141 77 143
rect 71 135 77 141
rect 58 134 77 135
rect 58 132 60 134
rect 62 132 77 134
rect 58 131 77 132
rect 55 120 56 122
rect 24 117 43 118
rect 24 115 39 117
rect 41 115 43 117
rect 24 114 43 115
rect 67 118 71 131
rect 98 139 99 145
rect 102 144 106 165
rect 125 147 129 165
rect 125 145 126 147
rect 128 145 129 147
rect 102 143 110 144
rect 102 141 106 143
rect 108 141 110 143
rect 102 140 110 141
rect 114 143 120 144
rect 125 143 129 145
rect 114 141 116 143
rect 118 141 120 143
rect 114 135 120 141
rect 101 134 120 135
rect 101 132 103 134
rect 105 132 120 134
rect 101 131 120 132
rect 98 120 99 122
rect 67 117 86 118
rect 67 115 82 117
rect 84 115 86 117
rect 67 114 86 115
rect 110 118 114 131
rect 141 139 142 145
rect 145 144 149 165
rect 168 147 172 165
rect 168 145 169 147
rect 171 145 172 147
rect 145 143 153 144
rect 145 141 149 143
rect 151 141 153 143
rect 145 140 153 141
rect 157 143 163 144
rect 168 143 172 145
rect 157 141 159 143
rect 161 141 163 143
rect 157 135 163 141
rect 144 134 163 135
rect 144 132 146 134
rect 148 132 163 134
rect 144 131 163 132
rect 141 120 142 122
rect 110 117 129 118
rect 110 115 125 117
rect 127 115 129 117
rect 110 114 129 115
rect 153 118 157 131
rect 153 117 172 118
rect 153 115 168 117
rect 170 115 172 117
rect 153 114 172 115
rect 18 67 20 69
rect 22 67 24 69
rect 18 66 24 67
rect 53 67 55 69
rect 57 67 59 69
rect 53 62 59 67
rect 75 67 77 69
rect 79 67 81 69
rect 53 60 55 62
rect 57 60 59 62
rect 53 59 59 60
rect 66 61 70 63
rect 66 59 67 61
rect 69 59 70 61
rect 75 62 81 67
rect 75 60 77 62
rect 79 60 81 62
rect 75 59 81 60
rect 119 67 121 69
rect 123 67 125 69
rect 119 62 125 67
rect 141 67 143 69
rect 145 67 147 69
rect 119 60 121 62
rect 123 60 125 62
rect 119 59 125 60
rect 130 61 134 63
rect 130 59 131 61
rect 133 59 134 61
rect 141 62 147 67
rect 176 67 178 69
rect 180 67 182 69
rect 176 66 182 67
rect 141 60 143 62
rect 145 60 147 62
rect 141 59 147 60
rect 23 55 47 59
rect 66 55 70 59
rect 21 51 27 55
rect 43 54 83 55
rect 43 52 67 54
rect 69 52 83 54
rect 21 41 25 51
rect 31 50 35 52
rect 43 51 83 52
rect 31 48 32 50
rect 34 48 35 50
rect 31 47 35 48
rect 21 39 22 41
rect 24 39 25 41
rect 21 37 25 39
rect 28 43 35 47
rect 28 32 32 43
rect 71 38 75 43
rect 71 36 72 38
rect 74 36 75 38
rect 71 34 75 36
rect 79 40 83 51
rect 79 38 85 40
rect 79 36 82 38
rect 84 36 85 38
rect 79 34 85 36
rect 14 31 32 32
rect 14 29 16 31
rect 18 30 32 31
rect 18 29 43 30
rect 14 28 39 29
rect 28 27 39 28
rect 41 27 43 29
rect 28 26 43 27
rect 48 29 52 31
rect 48 27 49 29
rect 51 27 52 29
rect 48 22 52 27
rect 79 31 83 34
rect 63 27 83 31
rect 63 23 67 27
rect 27 21 49 22
rect 18 18 22 20
rect 27 19 29 21
rect 31 20 49 21
rect 51 20 52 22
rect 31 19 52 20
rect 57 22 67 23
rect 57 20 59 22
rect 61 20 67 22
rect 57 19 67 20
rect 130 55 134 59
rect 153 55 177 59
rect 117 54 157 55
rect 117 52 131 54
rect 133 52 157 54
rect 117 51 157 52
rect 117 40 121 51
rect 165 50 169 52
rect 173 51 179 55
rect 165 48 166 50
rect 168 48 169 50
rect 165 47 169 48
rect 165 43 172 47
rect 115 38 121 40
rect 115 36 116 38
rect 118 36 121 38
rect 115 34 121 36
rect 125 38 129 43
rect 125 36 126 38
rect 128 36 129 38
rect 125 34 129 36
rect 117 31 121 34
rect 117 27 137 31
rect 133 23 137 27
rect 168 32 172 43
rect 175 41 179 51
rect 175 39 176 41
rect 178 39 179 41
rect 175 37 179 39
rect 168 31 186 32
rect 148 29 152 31
rect 168 30 182 31
rect 148 27 149 29
rect 151 27 152 29
rect 133 22 143 23
rect 133 20 139 22
rect 141 20 143 22
rect 133 19 143 20
rect 148 22 152 27
rect 157 29 182 30
rect 184 29 186 31
rect 157 27 159 29
rect 161 28 186 29
rect 161 27 172 28
rect 157 26 172 27
rect 148 20 149 22
rect 151 21 173 22
rect 151 20 169 21
rect 148 19 169 20
rect 171 19 173 21
rect 27 18 52 19
rect 148 18 173 19
rect 178 18 182 20
rect 18 16 19 18
rect 21 16 22 18
rect 178 16 179 18
rect 181 16 182 18
rect 18 13 22 16
rect 74 15 80 16
rect 74 13 76 15
rect 78 13 80 15
rect 120 15 126 16
rect 120 13 122 15
rect 124 13 126 15
rect 178 13 182 16
<< via1 >>
rect 9 125 11 127
rect 52 124 54 126
rect 95 124 97 126
rect 48 44 50 46
rect 56 32 58 34
rect 158 44 160 46
rect 109 33 111 35
rect 136 36 138 38
<< labels >>
rlabel alu1 69 105 69 105 6 vss
rlabel alu1 112 169 112 169 6 vdd
rlabel alu1 147 9 147 9 4 vss
rlabel alu1 147 73 147 73 4 vdd
rlabel polyct1 37 125 37 125 1 x1
rlabel polyct1 28 157 28 157 1 y1
rlabel polyct1 71 157 71 157 1 x1
rlabel polyct1 80 125 80 125 1 yo
rlabel polyct1 157 157 157 157 1 yo
rlabel polyct1 166 125 166 125 1 xo
rlabel polyct1 123 125 123 125 1 xo
rlabel alu1 89 49 89 49 1 p3
rlabel alu1 9 37 9 37 1 p2
rlabel alu1 139 132 139 132 1 p0
rlabel alu1 191 37 191 37 1 p1
<< end >>
