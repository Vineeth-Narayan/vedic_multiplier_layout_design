magic
tech scmos
timestamp 1636113200
<< ab >>
rect 10 39 137 77
rect 10 30 97 39
rect 100 30 137 39
rect 10 26 137 30
rect 10 24 97 26
rect 99 24 137 26
rect 10 5 137 24
rect 141 5 232 77
<< nwell >>
rect 8 37 232 82
<< pwell >>
rect 8 0 232 37
<< poly >>
rect 19 71 21 75
rect 42 68 44 73
rect 49 68 51 73
rect 67 71 69 75
rect 77 71 79 75
rect 87 71 89 75
rect 32 59 34 64
rect 19 33 21 46
rect 32 43 34 46
rect 121 71 123 75
rect 128 71 130 75
rect 148 71 150 75
rect 108 62 110 66
rect 25 41 34 43
rect 25 39 27 41
rect 29 39 31 41
rect 42 40 44 43
rect 49 40 51 43
rect 67 40 69 43
rect 77 40 79 43
rect 87 40 89 43
rect 108 41 110 50
rect 121 48 123 53
rect 118 46 124 48
rect 118 44 120 46
rect 122 44 124 46
rect 118 42 124 44
rect 25 37 31 39
rect 19 31 25 33
rect 19 29 21 31
rect 23 29 25 31
rect 19 27 25 29
rect 19 24 21 27
rect 29 24 31 37
rect 39 38 45 40
rect 39 36 41 38
rect 43 36 45 38
rect 39 34 45 36
rect 49 38 71 40
rect 49 36 60 38
rect 62 36 67 38
rect 69 36 71 38
rect 49 34 71 36
rect 75 38 81 40
rect 75 36 77 38
rect 79 36 81 38
rect 75 34 81 36
rect 85 38 91 40
rect 85 36 87 38
rect 89 36 91 38
rect 85 34 91 36
rect 108 39 114 41
rect 108 37 110 39
rect 112 37 114 39
rect 108 35 114 37
rect 39 31 41 34
rect 49 31 51 34
rect 69 31 71 34
rect 76 31 78 34
rect 19 7 21 11
rect 29 9 31 14
rect 39 12 41 17
rect 49 12 51 17
rect 87 25 89 34
rect 108 26 110 35
rect 118 26 120 42
rect 128 40 130 53
rect 171 68 173 73
rect 178 68 180 73
rect 196 71 198 75
rect 206 71 208 75
rect 216 71 218 75
rect 161 59 163 64
rect 128 38 134 40
rect 128 36 130 38
rect 132 36 134 38
rect 128 34 134 36
rect 128 26 130 34
rect 148 33 150 46
rect 161 43 163 46
rect 154 41 163 43
rect 154 39 156 41
rect 158 39 160 41
rect 171 40 173 43
rect 178 40 180 43
rect 196 40 198 43
rect 206 40 208 43
rect 216 40 218 43
rect 154 37 160 39
rect 148 31 154 33
rect 148 29 150 31
rect 152 29 154 31
rect 148 27 154 29
rect 148 24 150 27
rect 158 24 160 37
rect 168 38 174 40
rect 168 36 170 38
rect 172 36 174 38
rect 168 34 174 36
rect 178 38 200 40
rect 178 36 189 38
rect 191 36 196 38
rect 198 36 200 38
rect 178 34 200 36
rect 204 38 210 40
rect 204 36 206 38
rect 208 36 210 38
rect 204 34 210 36
rect 214 38 220 40
rect 214 36 216 38
rect 218 36 220 38
rect 214 34 220 36
rect 168 31 170 34
rect 178 31 180 34
rect 198 31 200 34
rect 205 31 207 34
rect 108 16 110 20
rect 118 16 120 20
rect 128 16 130 20
rect 69 7 71 11
rect 76 7 78 11
rect 87 7 89 11
rect 148 7 150 11
rect 158 9 160 14
rect 168 12 170 17
rect 178 12 180 17
rect 216 25 218 34
rect 198 7 200 11
rect 205 7 207 11
rect 216 7 218 11
<< ndif >>
rect 34 24 39 31
rect 12 22 19 24
rect 12 20 14 22
rect 16 20 19 22
rect 12 18 19 20
rect 14 11 19 18
rect 21 18 29 24
rect 21 16 24 18
rect 26 16 29 18
rect 21 14 29 16
rect 31 21 39 24
rect 31 19 34 21
rect 36 19 39 21
rect 31 17 39 19
rect 41 29 49 31
rect 41 27 44 29
rect 46 27 49 29
rect 41 17 49 27
rect 51 29 58 31
rect 51 27 54 29
rect 56 27 58 29
rect 51 22 58 27
rect 64 24 69 31
rect 51 20 54 22
rect 56 20 58 22
rect 51 17 58 20
rect 62 22 69 24
rect 62 20 64 22
rect 66 20 69 22
rect 62 18 69 20
rect 31 14 36 17
rect 21 11 26 14
rect 64 11 69 18
rect 71 11 76 31
rect 78 25 85 31
rect 78 15 87 25
rect 78 13 81 15
rect 83 13 87 15
rect 78 11 87 13
rect 89 22 96 25
rect 89 20 92 22
rect 94 20 96 22
rect 101 24 108 26
rect 101 22 103 24
rect 105 22 108 24
rect 101 20 108 22
rect 110 24 118 26
rect 110 22 113 24
rect 115 22 118 24
rect 110 20 118 22
rect 120 24 128 26
rect 120 22 123 24
rect 125 22 128 24
rect 120 20 128 22
rect 130 24 137 26
rect 163 24 168 31
rect 130 22 133 24
rect 135 22 137 24
rect 130 20 137 22
rect 141 22 148 24
rect 141 20 143 22
rect 145 20 148 22
rect 89 18 96 20
rect 89 11 94 18
rect 141 18 148 20
rect 143 11 148 18
rect 150 18 158 24
rect 150 16 153 18
rect 155 16 158 18
rect 150 14 158 16
rect 160 21 168 24
rect 160 19 163 21
rect 165 19 168 21
rect 160 17 168 19
rect 170 29 178 31
rect 170 27 173 29
rect 175 27 178 29
rect 170 17 178 27
rect 180 29 187 31
rect 180 27 183 29
rect 185 27 187 29
rect 180 22 187 27
rect 193 24 198 31
rect 180 20 183 22
rect 185 20 187 22
rect 180 17 187 20
rect 191 22 198 24
rect 191 20 193 22
rect 195 20 198 22
rect 191 18 198 20
rect 160 14 165 17
rect 150 11 155 14
rect 193 11 198 18
rect 200 11 205 31
rect 207 25 214 31
rect 207 15 216 25
rect 207 13 210 15
rect 212 13 216 15
rect 207 11 216 13
rect 218 22 225 25
rect 218 20 221 22
rect 223 20 225 22
rect 218 18 225 20
rect 218 11 223 18
<< pdif >>
rect 14 59 19 71
rect 12 57 19 59
rect 12 55 14 57
rect 16 55 19 57
rect 12 50 19 55
rect 12 48 14 50
rect 16 48 19 50
rect 12 46 19 48
rect 21 69 30 71
rect 21 67 25 69
rect 27 67 30 69
rect 53 69 67 71
rect 53 68 60 69
rect 21 59 30 67
rect 37 59 42 68
rect 21 46 32 59
rect 34 50 42 59
rect 34 48 37 50
rect 39 48 42 50
rect 34 46 42 48
rect 37 43 42 46
rect 44 43 49 68
rect 51 67 60 68
rect 62 67 67 69
rect 51 62 67 67
rect 51 60 60 62
rect 62 60 67 62
rect 51 43 67 60
rect 69 61 77 71
rect 69 59 72 61
rect 74 59 77 61
rect 69 54 77 59
rect 69 52 72 54
rect 74 52 77 54
rect 69 43 77 52
rect 79 69 87 71
rect 79 67 82 69
rect 84 67 87 69
rect 79 62 87 67
rect 79 60 82 62
rect 84 60 87 62
rect 79 43 87 60
rect 89 56 94 71
rect 112 69 121 71
rect 112 67 115 69
rect 117 67 121 69
rect 112 62 121 67
rect 101 60 108 62
rect 101 58 103 60
rect 105 58 108 60
rect 101 56 108 58
rect 89 54 96 56
rect 89 52 92 54
rect 94 52 96 54
rect 89 47 96 52
rect 103 50 108 56
rect 110 53 121 62
rect 123 53 128 71
rect 130 64 135 71
rect 130 62 137 64
rect 130 60 133 62
rect 135 60 137 62
rect 130 58 137 60
rect 143 59 148 71
rect 130 53 135 58
rect 141 57 148 59
rect 141 55 143 57
rect 145 55 148 57
rect 110 50 118 53
rect 89 45 92 47
rect 94 45 96 47
rect 89 43 96 45
rect 141 50 148 55
rect 141 48 143 50
rect 145 48 148 50
rect 141 46 148 48
rect 150 69 159 71
rect 150 67 154 69
rect 156 67 159 69
rect 182 69 196 71
rect 182 68 189 69
rect 150 59 159 67
rect 166 59 171 68
rect 150 46 161 59
rect 163 50 171 59
rect 163 48 166 50
rect 168 48 171 50
rect 163 46 171 48
rect 166 43 171 46
rect 173 43 178 68
rect 180 67 189 68
rect 191 67 196 69
rect 180 62 196 67
rect 180 60 189 62
rect 191 60 196 62
rect 180 43 196 60
rect 198 61 206 71
rect 198 59 201 61
rect 203 59 206 61
rect 198 54 206 59
rect 198 52 201 54
rect 203 52 206 54
rect 198 43 206 52
rect 208 69 216 71
rect 208 67 211 69
rect 213 67 216 69
rect 208 62 216 67
rect 208 60 211 62
rect 213 60 216 62
rect 208 43 216 60
rect 218 56 223 71
rect 218 54 225 56
rect 218 52 221 54
rect 223 52 225 54
rect 218 47 225 52
rect 218 45 221 47
rect 223 45 225 47
rect 218 43 225 45
<< alu1 >>
rect 8 72 232 77
rect 8 70 104 72
rect 106 70 232 72
rect 8 69 232 70
rect 12 59 25 63
rect 101 60 114 63
rect 12 57 17 59
rect 12 55 14 57
rect 16 55 17 57
rect 101 58 103 60
rect 105 59 114 60
rect 141 59 154 63
rect 12 50 17 55
rect 12 48 14 50
rect 16 48 17 50
rect 12 46 17 48
rect 12 24 16 46
rect 43 43 81 47
rect 43 40 48 43
rect 40 38 48 40
rect 40 36 41 38
rect 43 36 48 38
rect 40 34 48 36
rect 58 38 73 39
rect 58 36 60 38
rect 62 36 67 38
rect 69 36 73 38
rect 58 35 73 36
rect 12 22 17 24
rect 60 29 64 35
rect 91 54 97 56
rect 91 52 92 54
rect 94 52 97 54
rect 91 47 97 52
rect 91 45 92 47
rect 94 45 97 47
rect 91 43 97 45
rect 60 27 61 29
rect 63 27 64 29
rect 60 26 64 27
rect 93 23 97 43
rect 12 20 14 22
rect 16 20 17 22
rect 12 18 17 20
rect 75 22 97 23
rect 75 20 92 22
rect 94 20 97 22
rect 75 19 97 20
rect 101 26 105 58
rect 141 57 146 59
rect 125 47 129 56
rect 141 55 143 57
rect 145 55 146 57
rect 141 50 146 55
rect 141 48 143 50
rect 145 48 146 50
rect 116 46 129 47
rect 116 44 117 46
rect 119 44 120 46
rect 122 44 129 46
rect 116 43 129 44
rect 133 47 137 48
rect 133 45 134 47
rect 136 45 137 47
rect 133 39 137 45
rect 124 38 137 39
rect 124 36 130 38
rect 132 36 137 38
rect 124 35 137 36
rect 133 34 137 35
rect 141 46 146 48
rect 141 38 145 46
rect 141 36 142 38
rect 144 36 145 38
rect 172 43 210 47
rect 101 24 106 26
rect 101 22 103 24
rect 105 22 106 24
rect 101 18 106 22
rect 141 24 145 36
rect 172 40 177 43
rect 169 38 177 40
rect 169 36 170 38
rect 172 36 177 38
rect 169 34 177 36
rect 187 38 202 39
rect 187 36 189 38
rect 191 36 196 38
rect 198 36 202 38
rect 187 35 202 36
rect 141 22 146 24
rect 189 26 193 35
rect 220 54 226 56
rect 220 52 221 54
rect 223 52 226 54
rect 220 47 226 52
rect 220 45 221 47
rect 223 45 226 47
rect 220 43 226 45
rect 222 23 226 43
rect 141 20 143 22
rect 145 20 146 22
rect 141 18 146 20
rect 204 22 226 23
rect 204 20 221 22
rect 223 20 226 22
rect 204 19 226 20
rect 8 12 232 13
rect 8 10 104 12
rect 106 10 132 12
rect 134 10 232 12
rect 8 5 232 10
<< alu2 >>
rect 91 47 97 48
rect 133 47 224 48
rect 91 45 92 47
rect 94 46 120 47
rect 94 45 117 46
rect 91 44 117 45
rect 119 44 120 46
rect 133 45 134 47
rect 136 45 221 47
rect 223 45 224 47
rect 133 44 224 45
rect 91 43 120 44
rect 137 38 146 39
rect 137 36 142 38
rect 144 36 146 38
rect 137 35 146 36
rect 60 29 103 30
rect 137 29 141 35
rect 60 27 61 29
rect 63 27 141 29
rect 60 26 141 27
rect 99 24 141 26
<< ptie >>
rect 102 12 136 14
rect 102 10 104 12
rect 106 10 132 12
rect 134 10 136 12
rect 102 8 136 10
<< ntie >>
rect 102 72 108 74
rect 102 70 104 72
rect 106 70 108 72
rect 102 68 108 70
<< nmos >>
rect 19 11 21 24
rect 29 14 31 24
rect 39 17 41 31
rect 49 17 51 31
rect 69 11 71 31
rect 76 11 78 31
rect 87 11 89 25
rect 108 20 110 26
rect 118 20 120 26
rect 128 20 130 26
rect 148 11 150 24
rect 158 14 160 24
rect 168 17 170 31
rect 178 17 180 31
rect 198 11 200 31
rect 205 11 207 31
rect 216 11 218 25
<< pmos >>
rect 19 46 21 71
rect 32 46 34 59
rect 42 43 44 68
rect 49 43 51 68
rect 67 43 69 71
rect 77 43 79 71
rect 87 43 89 71
rect 108 50 110 62
rect 121 53 123 71
rect 128 53 130 71
rect 148 46 150 71
rect 161 46 163 59
rect 171 43 173 68
rect 178 43 180 68
rect 196 43 198 71
rect 206 43 208 71
rect 216 43 218 71
<< polyct0 >>
rect 27 39 29 41
rect 21 29 23 31
rect 77 36 79 38
rect 87 36 89 38
rect 110 37 112 39
rect 156 39 158 41
rect 150 29 152 31
rect 206 36 208 38
rect 216 36 218 38
<< polyct1 >>
rect 120 44 122 46
rect 41 36 43 38
rect 60 36 62 38
rect 67 36 69 38
rect 130 36 132 38
rect 170 36 172 38
rect 189 36 191 38
rect 196 36 198 38
<< ndifct0 >>
rect 24 16 26 18
rect 34 19 36 21
rect 44 27 46 29
rect 54 27 56 29
rect 54 20 56 22
rect 64 20 66 22
rect 81 13 83 15
rect 113 22 115 24
rect 123 22 125 24
rect 133 22 135 24
rect 153 16 155 18
rect 163 19 165 21
rect 173 27 175 29
rect 183 27 185 29
rect 183 20 185 22
rect 193 20 195 22
rect 210 13 212 15
<< ndifct1 >>
rect 14 20 16 22
rect 92 20 94 22
rect 103 22 105 24
rect 143 20 145 22
rect 221 20 223 22
<< ntiect1 >>
rect 104 70 106 72
<< ptiect1 >>
rect 104 10 106 12
rect 132 10 134 12
<< pdifct0 >>
rect 25 67 27 69
rect 37 48 39 50
rect 60 67 62 69
rect 60 60 62 62
rect 72 59 74 61
rect 72 52 74 54
rect 82 67 84 69
rect 82 60 84 62
rect 115 67 117 69
rect 133 60 135 62
rect 154 67 156 69
rect 166 48 168 50
rect 189 67 191 69
rect 189 60 191 62
rect 201 59 203 61
rect 201 52 203 54
rect 211 67 213 69
rect 211 60 213 62
<< pdifct1 >>
rect 14 55 16 57
rect 14 48 16 50
rect 103 58 105 60
rect 92 52 94 54
rect 143 55 145 57
rect 92 45 94 47
rect 143 48 145 50
rect 221 52 223 54
rect 221 45 223 47
<< alu0 >>
rect 23 67 25 69
rect 27 67 29 69
rect 23 66 29 67
rect 58 67 60 69
rect 62 67 64 69
rect 58 62 64 67
rect 80 67 82 69
rect 84 67 86 69
rect 58 60 60 62
rect 62 60 64 62
rect 58 59 64 60
rect 71 61 75 63
rect 71 59 72 61
rect 74 59 75 61
rect 80 62 86 67
rect 113 67 115 69
rect 117 67 119 69
rect 113 66 119 67
rect 152 67 154 69
rect 156 67 158 69
rect 152 66 158 67
rect 187 67 189 69
rect 191 67 193 69
rect 80 60 82 62
rect 84 60 86 62
rect 80 59 86 60
rect 28 55 52 59
rect 71 55 75 59
rect 117 62 137 63
rect 117 60 133 62
rect 135 60 137 62
rect 117 59 137 60
rect 187 62 193 67
rect 209 67 211 69
rect 213 67 215 69
rect 187 60 189 62
rect 191 60 193 62
rect 187 59 193 60
rect 200 61 204 63
rect 200 59 201 61
rect 203 59 204 61
rect 209 62 215 67
rect 209 60 211 62
rect 213 60 215 62
rect 209 59 215 60
rect 26 51 32 55
rect 48 54 88 55
rect 48 52 72 54
rect 74 52 88 54
rect 26 41 30 51
rect 36 50 40 52
rect 48 51 88 52
rect 36 48 37 50
rect 39 48 40 50
rect 36 47 40 48
rect 26 39 27 41
rect 29 39 30 41
rect 26 37 30 39
rect 33 43 40 47
rect 33 32 37 43
rect 76 38 80 43
rect 76 36 77 38
rect 79 36 80 38
rect 19 31 37 32
rect 19 29 21 31
rect 23 30 37 31
rect 23 29 48 30
rect 19 28 44 29
rect 33 27 44 28
rect 46 27 48 29
rect 33 26 48 27
rect 53 29 57 31
rect 53 27 54 29
rect 56 27 57 29
rect 53 22 57 27
rect 76 34 80 36
rect 84 40 88 51
rect 84 38 90 40
rect 84 36 87 38
rect 89 36 90 38
rect 84 34 90 36
rect 84 31 88 34
rect 68 27 88 31
rect 68 23 72 27
rect 32 21 54 22
rect 23 18 27 20
rect 32 19 34 21
rect 36 20 54 21
rect 56 20 57 22
rect 36 19 57 20
rect 62 22 72 23
rect 62 20 64 22
rect 66 20 72 22
rect 62 19 72 20
rect 105 56 106 59
rect 117 55 121 59
rect 109 51 121 55
rect 109 39 113 51
rect 157 55 181 59
rect 200 55 204 59
rect 109 37 110 39
rect 112 37 113 39
rect 109 32 113 37
rect 155 51 161 55
rect 177 54 217 55
rect 177 52 201 54
rect 203 52 217 54
rect 155 41 159 51
rect 165 50 169 52
rect 177 51 217 52
rect 165 48 166 50
rect 168 48 169 50
rect 165 47 169 48
rect 155 39 156 41
rect 158 39 159 41
rect 155 37 159 39
rect 162 43 169 47
rect 109 28 126 32
rect 32 18 57 19
rect 111 24 117 25
rect 111 22 113 24
rect 115 22 117 24
rect 23 16 24 18
rect 26 16 27 18
rect 23 13 27 16
rect 79 15 85 16
rect 79 13 81 15
rect 83 13 85 15
rect 111 13 117 22
rect 122 24 126 28
rect 122 22 123 24
rect 125 22 126 24
rect 122 20 126 22
rect 131 24 137 25
rect 131 22 133 24
rect 135 22 137 24
rect 131 13 137 22
rect 162 32 166 43
rect 205 38 209 43
rect 205 36 206 38
rect 208 36 209 38
rect 148 31 166 32
rect 148 29 150 31
rect 152 30 166 31
rect 152 29 177 30
rect 148 28 173 29
rect 162 27 173 28
rect 175 27 177 29
rect 162 26 177 27
rect 182 29 186 31
rect 182 27 183 29
rect 185 27 186 29
rect 182 22 186 27
rect 205 34 209 36
rect 213 40 217 51
rect 213 38 219 40
rect 213 36 216 38
rect 218 36 219 38
rect 213 34 219 36
rect 213 31 217 34
rect 197 27 217 31
rect 197 23 201 27
rect 161 21 183 22
rect 152 18 156 20
rect 161 19 163 21
rect 165 20 183 21
rect 185 20 186 22
rect 165 19 186 20
rect 191 22 201 23
rect 191 20 193 22
rect 195 20 201 22
rect 191 19 201 20
rect 161 18 186 19
rect 152 16 153 18
rect 155 16 156 18
rect 152 13 156 16
rect 208 15 214 16
rect 208 13 210 15
rect 212 13 214 15
<< via1 >>
rect 92 45 94 47
rect 61 27 63 29
rect 117 44 119 46
rect 134 45 136 47
rect 142 36 144 38
rect 221 45 223 47
<< labels >>
rlabel alu1 103 37 103 37 1 co
rlabel alu1 191 33 191 33 6 a
rlabel alu1 183 45 183 45 6 b
rlabel alu1 70 45 70 45 1 ci
rlabel alu1 58 73 58 73 6 vdd
rlabel alu1 58 9 58 9 6 vss
rlabel alu1 14 37 14 37 6 so
<< end >>
