magic
tech scmos
timestamp 1636532566
<< ab >>
rect 73 331 169 381
rect 173 343 300 381
rect 173 334 260 343
rect 263 334 300 343
rect 73 330 160 331
rect 173 330 300 334
rect 73 317 169 330
rect 173 328 260 330
rect 262 328 300 330
rect 173 317 300 328
rect 73 313 154 317
rect 174 313 300 317
rect 73 309 169 313
rect 173 309 300 313
rect 304 309 395 381
rect 397 343 524 381
rect 397 334 484 343
rect 487 334 524 343
rect 397 330 524 334
rect 397 328 484 330
rect 486 328 524 330
rect 397 309 524 328
rect 528 309 619 381
rect 622 309 718 381
rect 721 309 761 381
rect 770 309 810 381
rect 820 309 860 381
rect 73 215 113 287
rect 123 215 163 287
rect 194 216 234 288
rect 235 216 275 288
rect 323 215 363 287
rect 373 215 413 287
rect 417 215 457 287
rect 473 274 513 287
rect 473 268 498 274
rect 503 268 513 274
rect 473 215 513 268
rect 523 215 563 287
rect 573 274 613 287
rect 573 268 598 274
rect 603 268 613 274
rect 573 215 613 268
rect 623 215 663 287
rect 667 215 763 287
rect 767 215 863 287
rect 866 215 867 287
rect 73 155 200 193
rect 73 146 160 155
rect 163 146 200 155
rect 73 142 200 146
rect 73 140 160 142
rect 162 140 200 142
rect 73 121 200 140
rect 204 128 295 193
rect 204 121 232 128
rect 238 121 295 128
rect 297 155 424 193
rect 297 146 384 155
rect 387 146 424 155
rect 297 134 298 146
rect 303 142 424 146
rect 303 140 384 142
rect 386 140 424 142
rect 303 134 424 140
rect 297 121 424 134
rect 428 121 519 193
rect 521 155 648 193
rect 521 146 608 155
rect 611 146 648 155
rect 521 142 648 146
rect 521 140 608 142
rect 610 140 648 142
rect 521 121 648 140
rect 652 121 743 193
rect 745 121 785 193
rect 72 27 112 99
rect 116 61 243 99
rect 116 52 203 61
rect 206 52 243 61
rect 116 48 243 52
rect 116 46 203 48
rect 205 46 243 48
rect 116 36 243 46
rect 116 27 201 36
rect 217 27 243 36
rect 247 27 338 99
rect 339 27 379 99
rect 382 61 509 99
rect 382 52 469 61
rect 472 52 509 61
rect 382 48 509 52
rect 382 46 469 48
rect 471 46 509 48
rect 382 36 509 46
rect 382 27 464 36
rect 482 27 509 36
rect 513 27 604 99
rect 606 27 646 99
rect 648 61 775 99
rect 648 52 735 61
rect 738 52 775 61
rect 648 48 775 52
rect 648 46 735 48
rect 737 46 775 48
rect 648 41 775 46
rect 648 37 743 41
rect 744 37 775 41
rect 648 35 733 37
rect 648 27 732 35
rect 748 27 775 37
rect 779 27 870 99
rect 871 27 911 99
<< nwell >>
rect 68 341 865 386
rect 68 289 170 292
rect 314 289 457 292
rect 495 289 867 292
rect 68 248 867 289
rect 68 247 230 248
rect 165 245 230 247
rect 296 247 867 248
rect 296 245 316 247
rect 457 246 491 247
rect 82 195 590 198
rect 637 195 786 198
rect 82 193 786 195
rect 71 153 786 193
rect 67 99 524 104
rect 760 99 916 104
rect 67 59 916 99
<< pwell >>
rect 68 304 865 341
rect 68 245 165 247
rect 230 245 280 248
rect 316 246 457 247
rect 491 246 867 247
rect 316 245 867 246
rect 68 210 167 245
rect 189 211 280 245
rect 315 211 867 245
rect 315 210 786 211
rect 71 120 786 153
rect 71 119 505 120
rect 538 119 556 120
rect 71 117 316 119
rect 540 117 556 119
rect 71 116 294 117
rect 678 116 786 120
rect 67 22 916 59
rect 725 14 821 22
rect 725 8 766 14
<< poly >>
rect 82 375 84 379
rect 105 372 107 377
rect 112 372 114 377
rect 130 375 132 379
rect 140 375 142 379
rect 150 375 152 379
rect 182 375 184 379
rect 95 363 97 368
rect 82 337 84 350
rect 95 347 97 350
rect 205 372 207 377
rect 212 372 214 377
rect 230 375 232 379
rect 240 375 242 379
rect 250 375 252 379
rect 195 363 197 368
rect 88 345 97 347
rect 88 343 90 345
rect 92 343 94 345
rect 105 344 107 347
rect 112 344 114 347
rect 130 344 132 347
rect 140 344 142 347
rect 150 344 152 347
rect 88 341 94 343
rect 82 335 88 337
rect 82 333 84 335
rect 86 333 88 335
rect 82 331 88 333
rect 82 328 84 331
rect 92 328 94 341
rect 102 342 108 344
rect 102 340 104 342
rect 106 340 108 342
rect 102 338 108 340
rect 112 342 134 344
rect 112 340 123 342
rect 125 340 130 342
rect 132 340 134 342
rect 112 338 134 340
rect 138 342 144 344
rect 138 340 140 342
rect 142 340 144 342
rect 138 338 144 340
rect 148 342 154 344
rect 148 340 150 342
rect 152 340 154 342
rect 148 338 154 340
rect 102 335 104 338
rect 112 335 114 338
rect 132 335 134 338
rect 139 335 141 338
rect 82 311 84 315
rect 92 313 94 318
rect 102 316 104 321
rect 112 316 114 321
rect 150 329 152 338
rect 182 337 184 350
rect 195 347 197 350
rect 284 375 286 379
rect 291 375 293 379
rect 311 375 313 379
rect 271 366 273 370
rect 188 345 197 347
rect 188 343 190 345
rect 192 343 194 345
rect 205 344 207 347
rect 212 344 214 347
rect 230 344 232 347
rect 240 344 242 347
rect 250 344 252 347
rect 271 345 273 354
rect 284 352 286 357
rect 281 350 287 352
rect 281 348 283 350
rect 285 348 287 350
rect 281 346 287 348
rect 188 341 194 343
rect 182 335 188 337
rect 182 333 184 335
rect 186 333 188 335
rect 182 331 188 333
rect 182 328 184 331
rect 192 328 194 341
rect 202 342 208 344
rect 202 340 204 342
rect 206 340 208 342
rect 202 338 208 340
rect 212 342 234 344
rect 212 340 223 342
rect 225 340 230 342
rect 232 340 234 342
rect 212 338 234 340
rect 238 342 244 344
rect 238 340 240 342
rect 242 340 244 342
rect 238 338 244 340
rect 248 342 254 344
rect 248 340 250 342
rect 252 340 254 342
rect 248 338 254 340
rect 271 343 277 345
rect 271 341 273 343
rect 275 341 277 343
rect 271 339 277 341
rect 202 335 204 338
rect 212 335 214 338
rect 232 335 234 338
rect 239 335 241 338
rect 132 311 134 315
rect 139 311 141 315
rect 150 311 152 315
rect 182 311 184 315
rect 192 313 194 318
rect 202 316 204 321
rect 212 316 214 321
rect 250 329 252 338
rect 271 330 273 339
rect 281 330 283 346
rect 291 344 293 357
rect 334 372 336 377
rect 341 372 343 377
rect 359 375 361 379
rect 369 375 371 379
rect 379 375 381 379
rect 406 375 408 379
rect 324 363 326 368
rect 291 342 297 344
rect 291 340 293 342
rect 295 340 297 342
rect 291 338 297 340
rect 291 330 293 338
rect 311 337 313 350
rect 324 347 326 350
rect 429 372 431 377
rect 436 372 438 377
rect 454 375 456 379
rect 464 375 466 379
rect 474 375 476 379
rect 419 363 421 368
rect 317 345 326 347
rect 317 343 319 345
rect 321 343 323 345
rect 334 344 336 347
rect 341 344 343 347
rect 359 344 361 347
rect 369 344 371 347
rect 379 344 381 347
rect 317 341 323 343
rect 311 335 317 337
rect 311 333 313 335
rect 315 333 317 335
rect 311 331 317 333
rect 311 328 313 331
rect 321 328 323 341
rect 331 342 337 344
rect 331 340 333 342
rect 335 340 337 342
rect 331 338 337 340
rect 341 342 363 344
rect 341 340 352 342
rect 354 340 359 342
rect 361 340 363 342
rect 341 338 363 340
rect 367 342 373 344
rect 367 340 369 342
rect 371 340 373 342
rect 367 338 373 340
rect 377 342 383 344
rect 377 340 379 342
rect 381 340 383 342
rect 377 338 383 340
rect 331 335 333 338
rect 341 335 343 338
rect 361 335 363 338
rect 368 335 370 338
rect 271 320 273 324
rect 281 320 283 324
rect 291 320 293 324
rect 232 311 234 315
rect 239 311 241 315
rect 250 311 252 315
rect 311 311 313 315
rect 321 313 323 318
rect 331 316 333 321
rect 341 316 343 321
rect 379 329 381 338
rect 406 337 408 350
rect 419 347 421 350
rect 508 375 510 379
rect 515 375 517 379
rect 535 375 537 379
rect 495 366 497 370
rect 412 345 421 347
rect 412 343 414 345
rect 416 343 418 345
rect 429 344 431 347
rect 436 344 438 347
rect 454 344 456 347
rect 464 344 466 347
rect 474 344 476 347
rect 495 345 497 354
rect 508 352 510 357
rect 505 350 511 352
rect 505 348 507 350
rect 509 348 511 350
rect 505 346 511 348
rect 412 341 418 343
rect 406 335 412 337
rect 406 333 408 335
rect 410 333 412 335
rect 406 331 412 333
rect 406 328 408 331
rect 416 328 418 341
rect 426 342 432 344
rect 426 340 428 342
rect 430 340 432 342
rect 426 338 432 340
rect 436 342 458 344
rect 436 340 447 342
rect 449 340 454 342
rect 456 340 458 342
rect 436 338 458 340
rect 462 342 468 344
rect 462 340 464 342
rect 466 340 468 342
rect 462 338 468 340
rect 472 342 478 344
rect 472 340 474 342
rect 476 340 478 342
rect 472 338 478 340
rect 495 343 501 345
rect 495 341 497 343
rect 499 341 501 343
rect 495 339 501 341
rect 426 335 428 338
rect 436 335 438 338
rect 456 335 458 338
rect 463 335 465 338
rect 361 311 363 315
rect 368 311 370 315
rect 379 311 381 315
rect 406 311 408 315
rect 416 313 418 318
rect 426 316 428 321
rect 436 316 438 321
rect 474 329 476 338
rect 495 330 497 339
rect 505 330 507 346
rect 515 344 517 357
rect 558 372 560 377
rect 565 372 567 377
rect 583 375 585 379
rect 593 375 595 379
rect 603 375 605 379
rect 631 375 633 379
rect 548 363 550 368
rect 515 342 521 344
rect 515 340 517 342
rect 519 340 521 342
rect 515 338 521 340
rect 515 330 517 338
rect 535 337 537 350
rect 548 347 550 350
rect 654 372 656 377
rect 661 372 663 377
rect 679 375 681 379
rect 689 375 691 379
rect 699 375 701 379
rect 644 363 646 368
rect 541 345 550 347
rect 541 343 543 345
rect 545 343 547 345
rect 558 344 560 347
rect 565 344 567 347
rect 583 344 585 347
rect 593 344 595 347
rect 603 344 605 347
rect 541 341 547 343
rect 535 335 541 337
rect 535 333 537 335
rect 539 333 541 335
rect 535 331 541 333
rect 535 328 537 331
rect 545 328 547 341
rect 555 342 561 344
rect 555 340 557 342
rect 559 340 561 342
rect 555 338 561 340
rect 565 342 587 344
rect 565 340 576 342
rect 578 340 583 342
rect 585 340 587 342
rect 565 338 587 340
rect 591 342 597 344
rect 591 340 593 342
rect 595 340 597 342
rect 591 338 597 340
rect 601 342 607 344
rect 601 340 603 342
rect 605 340 607 342
rect 601 338 607 340
rect 555 335 557 338
rect 565 335 567 338
rect 585 335 587 338
rect 592 335 594 338
rect 495 320 497 324
rect 505 320 507 324
rect 515 320 517 324
rect 456 311 458 315
rect 463 311 465 315
rect 474 311 476 315
rect 535 311 537 315
rect 545 313 547 318
rect 555 316 557 321
rect 565 316 567 321
rect 603 329 605 338
rect 631 337 633 350
rect 644 347 646 350
rect 740 366 746 368
rect 740 364 742 366
rect 744 364 746 366
rect 789 366 795 368
rect 789 364 791 366
rect 793 364 795 366
rect 839 366 845 368
rect 839 364 841 366
rect 843 364 845 366
rect 730 359 732 364
rect 740 362 746 364
rect 740 357 742 362
rect 750 357 752 362
rect 779 359 781 364
rect 789 362 795 364
rect 789 357 791 362
rect 799 357 801 362
rect 829 359 831 364
rect 839 362 845 364
rect 839 357 841 362
rect 849 357 851 362
rect 637 345 646 347
rect 637 343 639 345
rect 641 343 643 345
rect 654 344 656 347
rect 661 344 663 347
rect 679 344 681 347
rect 689 344 691 347
rect 699 344 701 347
rect 730 344 732 347
rect 740 344 742 347
rect 637 341 643 343
rect 631 335 637 337
rect 631 333 633 335
rect 635 333 637 335
rect 631 331 637 333
rect 631 328 633 331
rect 641 328 643 341
rect 651 342 657 344
rect 651 340 653 342
rect 655 340 657 342
rect 651 338 657 340
rect 661 342 683 344
rect 661 340 672 342
rect 674 340 679 342
rect 681 340 683 342
rect 661 338 683 340
rect 687 342 693 344
rect 687 340 689 342
rect 691 340 693 342
rect 687 338 693 340
rect 697 342 703 344
rect 697 340 699 342
rect 701 340 703 342
rect 697 338 703 340
rect 730 342 736 344
rect 730 340 732 342
rect 734 340 736 342
rect 740 341 744 344
rect 730 338 736 340
rect 651 335 653 338
rect 661 335 663 338
rect 681 335 683 338
rect 688 335 690 338
rect 585 311 587 315
rect 592 311 594 315
rect 603 311 605 315
rect 631 311 633 315
rect 641 313 643 318
rect 651 316 653 321
rect 661 316 663 321
rect 699 329 701 338
rect 730 330 732 338
rect 742 327 744 341
rect 750 336 752 347
rect 779 344 781 347
rect 789 344 791 347
rect 779 342 785 344
rect 779 340 781 342
rect 783 340 785 342
rect 789 341 793 344
rect 779 338 785 340
rect 749 334 755 336
rect 749 332 751 334
rect 753 332 755 334
rect 749 330 755 332
rect 779 330 781 338
rect 749 327 751 330
rect 730 320 732 324
rect 791 327 793 341
rect 799 336 801 347
rect 829 344 831 347
rect 839 344 841 347
rect 829 342 835 344
rect 829 340 831 342
rect 833 340 835 342
rect 839 341 843 344
rect 829 338 835 340
rect 798 334 804 336
rect 798 332 800 334
rect 802 332 804 334
rect 798 330 804 332
rect 829 330 831 338
rect 798 327 800 330
rect 779 320 781 324
rect 841 327 843 341
rect 849 336 851 347
rect 848 334 854 336
rect 848 332 850 334
rect 852 332 854 334
rect 848 330 854 332
rect 848 327 850 330
rect 829 320 831 324
rect 681 311 683 315
rect 688 311 690 315
rect 699 311 701 315
rect 742 313 744 318
rect 749 313 751 318
rect 791 313 793 318
rect 798 313 800 318
rect 841 313 843 318
rect 848 313 850 318
rect 676 281 678 285
rect 92 272 98 274
rect 92 270 94 272
rect 96 270 98 272
rect 142 272 148 274
rect 142 270 144 272
rect 146 270 148 272
rect 213 273 219 275
rect 213 271 215 273
rect 217 271 219 273
rect 254 273 260 275
rect 254 271 256 273
rect 258 271 260 273
rect 82 265 84 270
rect 92 268 98 270
rect 92 263 94 268
rect 102 263 104 268
rect 132 265 134 270
rect 142 268 148 270
rect 142 263 144 268
rect 152 263 154 268
rect 203 266 205 271
rect 213 269 219 271
rect 213 264 215 269
rect 223 264 225 269
rect 244 266 246 271
rect 254 269 260 271
rect 342 272 348 274
rect 342 270 344 272
rect 346 270 348 272
rect 392 272 398 274
rect 392 270 394 272
rect 396 270 398 272
rect 436 272 442 274
rect 436 270 438 272
rect 440 270 442 272
rect 492 272 498 274
rect 492 270 494 272
rect 496 270 498 272
rect 542 272 548 274
rect 542 270 544 272
rect 546 270 548 272
rect 592 272 598 274
rect 592 270 594 272
rect 596 270 598 272
rect 642 272 648 274
rect 642 270 644 272
rect 646 270 648 272
rect 254 264 256 269
rect 264 264 266 269
rect 332 265 334 270
rect 342 268 348 270
rect 82 250 84 253
rect 92 250 94 253
rect 82 248 88 250
rect 82 246 84 248
rect 86 246 88 248
rect 92 247 96 250
rect 82 244 88 246
rect 82 236 84 244
rect 94 233 96 247
rect 102 242 104 253
rect 132 250 134 253
rect 142 250 144 253
rect 132 248 138 250
rect 132 246 134 248
rect 136 246 138 248
rect 142 247 146 250
rect 132 244 138 246
rect 101 240 107 242
rect 101 238 103 240
rect 105 238 107 240
rect 101 236 107 238
rect 132 236 134 244
rect 101 233 103 236
rect 82 226 84 230
rect 144 233 146 247
rect 152 242 154 253
rect 203 251 205 254
rect 213 251 215 254
rect 203 249 209 251
rect 203 247 205 249
rect 207 247 209 249
rect 213 248 217 251
rect 203 245 209 247
rect 151 240 157 242
rect 151 238 153 240
rect 155 238 157 240
rect 151 236 157 238
rect 203 237 205 245
rect 151 233 153 236
rect 132 226 134 230
rect 215 234 217 248
rect 223 243 225 254
rect 244 251 246 254
rect 254 251 256 254
rect 244 249 250 251
rect 244 247 246 249
rect 248 247 250 249
rect 254 248 258 251
rect 244 245 250 247
rect 222 241 228 243
rect 222 239 224 241
rect 226 239 228 241
rect 222 237 228 239
rect 244 237 246 245
rect 222 234 224 237
rect 203 227 205 231
rect 256 234 258 248
rect 264 243 266 254
rect 342 263 344 268
rect 352 263 354 268
rect 382 265 384 270
rect 392 268 398 270
rect 392 263 394 268
rect 402 263 404 268
rect 426 265 428 270
rect 436 268 442 270
rect 436 263 438 268
rect 446 263 448 268
rect 482 265 484 270
rect 492 268 498 270
rect 492 263 494 268
rect 502 263 504 268
rect 532 265 534 270
rect 542 268 548 270
rect 542 263 544 268
rect 552 263 554 268
rect 582 265 584 270
rect 592 268 598 270
rect 592 263 594 268
rect 602 263 604 268
rect 632 265 634 270
rect 642 268 648 270
rect 642 263 644 268
rect 652 263 654 268
rect 699 278 701 283
rect 706 278 708 283
rect 724 281 726 285
rect 734 281 736 285
rect 744 281 746 285
rect 776 281 778 285
rect 689 269 691 274
rect 332 250 334 253
rect 342 250 344 253
rect 332 248 338 250
rect 332 246 334 248
rect 336 246 338 248
rect 342 247 346 250
rect 332 244 338 246
rect 263 241 269 243
rect 263 239 265 241
rect 267 239 269 241
rect 263 237 269 239
rect 263 234 265 237
rect 332 236 334 244
rect 244 227 246 231
rect 344 233 346 247
rect 352 242 354 253
rect 382 250 384 253
rect 392 250 394 253
rect 382 248 388 250
rect 382 246 384 248
rect 386 246 388 248
rect 392 247 396 250
rect 382 244 388 246
rect 351 240 357 242
rect 351 238 353 240
rect 355 238 357 240
rect 351 236 357 238
rect 382 236 384 244
rect 351 233 353 236
rect 332 226 334 230
rect 94 219 96 224
rect 101 219 103 224
rect 144 219 146 224
rect 151 219 153 224
rect 215 220 217 225
rect 222 220 224 225
rect 256 220 258 225
rect 263 220 265 225
rect 394 233 396 247
rect 402 242 404 253
rect 426 250 428 253
rect 436 250 438 253
rect 426 248 432 250
rect 426 246 428 248
rect 430 246 432 248
rect 436 247 440 250
rect 426 244 432 246
rect 401 240 407 242
rect 401 238 403 240
rect 405 238 407 240
rect 401 236 407 238
rect 426 236 428 244
rect 401 233 403 236
rect 382 226 384 230
rect 438 233 440 247
rect 446 242 448 253
rect 482 250 484 253
rect 492 250 494 253
rect 482 248 488 250
rect 482 246 484 248
rect 486 246 488 248
rect 492 247 496 250
rect 482 244 488 246
rect 445 240 451 242
rect 445 238 447 240
rect 449 238 451 240
rect 445 236 451 238
rect 482 236 484 244
rect 445 233 447 236
rect 426 226 428 230
rect 494 233 496 247
rect 502 242 504 253
rect 532 250 534 253
rect 542 250 544 253
rect 532 248 538 250
rect 532 246 534 248
rect 536 246 538 248
rect 542 247 546 250
rect 532 244 538 246
rect 501 240 507 242
rect 501 238 503 240
rect 505 238 507 240
rect 501 236 507 238
rect 532 236 534 244
rect 501 233 503 236
rect 482 226 484 230
rect 544 233 546 247
rect 552 242 554 253
rect 582 250 584 253
rect 592 250 594 253
rect 582 248 588 250
rect 582 246 584 248
rect 586 246 588 248
rect 592 247 596 250
rect 582 244 588 246
rect 551 240 557 242
rect 551 238 553 240
rect 555 238 557 240
rect 551 236 557 238
rect 582 236 584 244
rect 551 233 553 236
rect 532 226 534 230
rect 594 233 596 247
rect 602 242 604 253
rect 632 250 634 253
rect 642 250 644 253
rect 632 248 638 250
rect 632 246 634 248
rect 636 246 638 248
rect 642 247 646 250
rect 632 244 638 246
rect 601 240 607 242
rect 601 238 603 240
rect 605 238 607 240
rect 601 236 607 238
rect 632 236 634 244
rect 601 233 603 236
rect 582 226 584 230
rect 644 233 646 247
rect 652 242 654 253
rect 676 243 678 256
rect 689 253 691 256
rect 799 278 801 283
rect 806 278 808 283
rect 824 281 826 285
rect 834 281 836 285
rect 844 281 846 285
rect 789 269 791 274
rect 682 251 691 253
rect 682 249 684 251
rect 686 249 688 251
rect 699 250 701 253
rect 706 250 708 253
rect 724 250 726 253
rect 734 250 736 253
rect 744 250 746 253
rect 682 247 688 249
rect 651 240 657 242
rect 651 238 653 240
rect 655 238 657 240
rect 651 236 657 238
rect 676 241 682 243
rect 676 239 678 241
rect 680 239 682 241
rect 676 237 682 239
rect 651 233 653 236
rect 676 234 678 237
rect 686 234 688 247
rect 696 248 702 250
rect 696 246 698 248
rect 700 246 702 248
rect 696 244 702 246
rect 706 248 728 250
rect 706 246 717 248
rect 719 246 724 248
rect 726 246 728 248
rect 706 244 728 246
rect 732 248 738 250
rect 732 246 734 248
rect 736 246 738 248
rect 732 244 738 246
rect 742 248 748 250
rect 742 246 744 248
rect 746 246 748 248
rect 742 244 748 246
rect 696 241 698 244
rect 706 241 708 244
rect 726 241 728 244
rect 733 241 735 244
rect 632 226 634 230
rect 344 219 346 224
rect 351 219 353 224
rect 394 219 396 224
rect 401 219 403 224
rect 438 219 440 224
rect 445 219 447 224
rect 494 219 496 224
rect 501 219 503 224
rect 544 219 546 224
rect 551 219 553 224
rect 594 219 596 224
rect 601 219 603 224
rect 644 219 646 224
rect 651 219 653 224
rect 676 217 678 221
rect 686 219 688 224
rect 696 222 698 227
rect 706 222 708 227
rect 744 235 746 244
rect 776 243 778 256
rect 789 253 791 256
rect 782 251 791 253
rect 782 249 784 251
rect 786 249 788 251
rect 799 250 801 253
rect 806 250 808 253
rect 824 250 826 253
rect 834 250 836 253
rect 844 250 846 253
rect 782 247 788 249
rect 776 241 782 243
rect 776 239 778 241
rect 780 239 782 241
rect 776 237 782 239
rect 776 234 778 237
rect 786 234 788 247
rect 796 248 802 250
rect 796 246 798 248
rect 800 246 802 248
rect 796 244 802 246
rect 806 248 828 250
rect 806 246 817 248
rect 819 246 824 248
rect 826 246 828 248
rect 806 244 828 246
rect 832 248 838 250
rect 832 246 834 248
rect 836 246 838 248
rect 832 244 838 246
rect 842 248 848 250
rect 842 246 844 248
rect 846 246 848 248
rect 842 244 848 246
rect 796 241 798 244
rect 806 241 808 244
rect 826 241 828 244
rect 833 241 835 244
rect 726 217 728 221
rect 733 217 735 221
rect 744 217 746 221
rect 776 217 778 221
rect 786 219 788 224
rect 796 222 798 227
rect 806 222 808 227
rect 844 235 846 244
rect 826 217 828 221
rect 833 217 835 221
rect 844 217 846 221
rect 82 187 84 191
rect 105 184 107 189
rect 112 184 114 189
rect 130 187 132 191
rect 140 187 142 191
rect 150 187 152 191
rect 95 175 97 180
rect 82 149 84 162
rect 95 159 97 162
rect 184 187 186 191
rect 191 187 193 191
rect 211 187 213 191
rect 171 178 173 182
rect 88 157 97 159
rect 88 155 90 157
rect 92 155 94 157
rect 105 156 107 159
rect 112 156 114 159
rect 130 156 132 159
rect 140 156 142 159
rect 150 156 152 159
rect 171 157 173 166
rect 184 164 186 169
rect 181 162 187 164
rect 181 160 183 162
rect 185 160 187 162
rect 181 158 187 160
rect 88 153 94 155
rect 82 147 88 149
rect 82 145 84 147
rect 86 145 88 147
rect 82 143 88 145
rect 82 140 84 143
rect 92 140 94 153
rect 102 154 108 156
rect 102 152 104 154
rect 106 152 108 154
rect 102 150 108 152
rect 112 154 134 156
rect 112 152 123 154
rect 125 152 130 154
rect 132 152 134 154
rect 112 150 134 152
rect 138 154 144 156
rect 138 152 140 154
rect 142 152 144 154
rect 138 150 144 152
rect 148 154 154 156
rect 148 152 150 154
rect 152 152 154 154
rect 148 150 154 152
rect 171 155 177 157
rect 171 153 173 155
rect 175 153 177 155
rect 171 151 177 153
rect 102 147 104 150
rect 112 147 114 150
rect 132 147 134 150
rect 139 147 141 150
rect 82 123 84 127
rect 92 125 94 130
rect 102 128 104 133
rect 112 128 114 133
rect 150 141 152 150
rect 171 142 173 151
rect 181 142 183 158
rect 191 156 193 169
rect 234 184 236 189
rect 241 184 243 189
rect 259 187 261 191
rect 269 187 271 191
rect 279 187 281 191
rect 306 187 308 191
rect 224 175 226 180
rect 191 154 197 156
rect 191 152 193 154
rect 195 152 197 154
rect 191 150 197 152
rect 191 142 193 150
rect 211 149 213 162
rect 224 159 226 162
rect 329 184 331 189
rect 336 184 338 189
rect 354 187 356 191
rect 364 187 366 191
rect 374 187 376 191
rect 319 175 321 180
rect 217 157 226 159
rect 217 155 219 157
rect 221 155 223 157
rect 234 156 236 159
rect 241 156 243 159
rect 259 156 261 159
rect 269 156 271 159
rect 279 156 281 159
rect 217 153 223 155
rect 211 147 217 149
rect 211 145 213 147
rect 215 145 217 147
rect 211 143 217 145
rect 211 140 213 143
rect 221 140 223 153
rect 231 154 237 156
rect 231 152 233 154
rect 235 152 237 154
rect 231 150 237 152
rect 241 154 263 156
rect 241 152 252 154
rect 254 152 259 154
rect 261 152 263 154
rect 241 150 263 152
rect 267 154 273 156
rect 267 152 269 154
rect 271 152 273 154
rect 267 150 273 152
rect 277 154 283 156
rect 277 152 279 154
rect 281 152 283 154
rect 277 150 283 152
rect 231 147 233 150
rect 241 147 243 150
rect 261 147 263 150
rect 268 147 270 150
rect 171 132 173 136
rect 181 132 183 136
rect 191 132 193 136
rect 132 123 134 127
rect 139 123 141 127
rect 150 123 152 127
rect 211 123 213 127
rect 221 125 223 130
rect 231 128 233 133
rect 241 128 243 133
rect 279 141 281 150
rect 306 149 308 162
rect 319 159 321 162
rect 408 187 410 191
rect 415 187 417 191
rect 435 187 437 191
rect 395 178 397 182
rect 312 157 321 159
rect 312 155 314 157
rect 316 155 318 157
rect 329 156 331 159
rect 336 156 338 159
rect 354 156 356 159
rect 364 156 366 159
rect 374 156 376 159
rect 395 157 397 166
rect 408 164 410 169
rect 405 162 411 164
rect 405 160 407 162
rect 409 160 411 162
rect 405 158 411 160
rect 312 153 318 155
rect 306 147 312 149
rect 306 145 308 147
rect 310 145 312 147
rect 306 143 312 145
rect 306 140 308 143
rect 316 140 318 153
rect 326 154 332 156
rect 326 152 328 154
rect 330 152 332 154
rect 326 150 332 152
rect 336 154 358 156
rect 336 152 347 154
rect 349 152 354 154
rect 356 152 358 154
rect 336 150 358 152
rect 362 154 368 156
rect 362 152 364 154
rect 366 152 368 154
rect 362 150 368 152
rect 372 154 378 156
rect 372 152 374 154
rect 376 152 378 154
rect 372 150 378 152
rect 395 155 401 157
rect 395 153 397 155
rect 399 153 401 155
rect 395 151 401 153
rect 326 147 328 150
rect 336 147 338 150
rect 356 147 358 150
rect 363 147 365 150
rect 261 123 263 127
rect 268 123 270 127
rect 279 123 281 127
rect 306 123 308 127
rect 316 125 318 130
rect 326 128 328 133
rect 336 128 338 133
rect 374 141 376 150
rect 395 142 397 151
rect 405 142 407 158
rect 415 156 417 169
rect 458 184 460 189
rect 465 184 467 189
rect 483 187 485 191
rect 493 187 495 191
rect 503 187 505 191
rect 530 187 532 191
rect 448 175 450 180
rect 415 154 421 156
rect 415 152 417 154
rect 419 152 421 154
rect 415 150 421 152
rect 415 142 417 150
rect 435 149 437 162
rect 448 159 450 162
rect 553 184 555 189
rect 560 184 562 189
rect 578 187 580 191
rect 588 187 590 191
rect 598 187 600 191
rect 543 175 545 180
rect 441 157 450 159
rect 441 155 443 157
rect 445 155 447 157
rect 458 156 460 159
rect 465 156 467 159
rect 483 156 485 159
rect 493 156 495 159
rect 503 156 505 159
rect 441 153 447 155
rect 435 147 441 149
rect 435 145 437 147
rect 439 145 441 147
rect 435 143 441 145
rect 435 140 437 143
rect 445 140 447 153
rect 455 154 461 156
rect 455 152 457 154
rect 459 152 461 154
rect 455 150 461 152
rect 465 154 487 156
rect 465 152 476 154
rect 478 152 483 154
rect 485 152 487 154
rect 465 150 487 152
rect 491 154 497 156
rect 491 152 493 154
rect 495 152 497 154
rect 491 150 497 152
rect 501 154 507 156
rect 501 152 503 154
rect 505 152 507 154
rect 501 150 507 152
rect 455 147 457 150
rect 465 147 467 150
rect 485 147 487 150
rect 492 147 494 150
rect 395 132 397 136
rect 405 132 407 136
rect 415 132 417 136
rect 356 123 358 127
rect 363 123 365 127
rect 374 123 376 127
rect 435 123 437 127
rect 445 125 447 130
rect 455 128 457 133
rect 465 128 467 133
rect 503 141 505 150
rect 530 149 532 162
rect 543 159 545 162
rect 632 187 634 191
rect 639 187 641 191
rect 659 187 661 191
rect 619 178 621 182
rect 536 157 545 159
rect 536 155 538 157
rect 540 155 542 157
rect 553 156 555 159
rect 560 156 562 159
rect 578 156 580 159
rect 588 156 590 159
rect 598 156 600 159
rect 619 157 621 166
rect 632 164 634 169
rect 629 162 635 164
rect 629 160 631 162
rect 633 160 635 162
rect 629 158 635 160
rect 536 153 542 155
rect 530 147 536 149
rect 530 145 532 147
rect 534 145 536 147
rect 530 143 536 145
rect 530 140 532 143
rect 540 140 542 153
rect 550 154 556 156
rect 550 152 552 154
rect 554 152 556 154
rect 550 150 556 152
rect 560 154 582 156
rect 560 152 571 154
rect 573 152 578 154
rect 580 152 582 154
rect 560 150 582 152
rect 586 154 592 156
rect 586 152 588 154
rect 590 152 592 154
rect 586 150 592 152
rect 596 154 602 156
rect 596 152 598 154
rect 600 152 602 154
rect 596 150 602 152
rect 619 155 625 157
rect 619 153 621 155
rect 623 153 625 155
rect 619 151 625 153
rect 550 147 552 150
rect 560 147 562 150
rect 580 147 582 150
rect 587 147 589 150
rect 485 123 487 127
rect 492 123 494 127
rect 503 123 505 127
rect 530 123 532 127
rect 540 125 542 130
rect 550 128 552 133
rect 560 128 562 133
rect 598 141 600 150
rect 619 142 621 151
rect 629 142 631 158
rect 639 156 641 169
rect 682 184 684 189
rect 689 184 691 189
rect 707 187 709 191
rect 717 187 719 191
rect 727 187 729 191
rect 672 175 674 180
rect 639 154 645 156
rect 639 152 641 154
rect 643 152 645 154
rect 639 150 645 152
rect 639 142 641 150
rect 659 149 661 162
rect 672 159 674 162
rect 764 178 770 180
rect 764 176 766 178
rect 768 176 770 178
rect 754 171 756 176
rect 764 174 770 176
rect 764 169 766 174
rect 774 169 776 174
rect 665 157 674 159
rect 665 155 667 157
rect 669 155 671 157
rect 682 156 684 159
rect 689 156 691 159
rect 707 156 709 159
rect 717 156 719 159
rect 727 156 729 159
rect 754 156 756 159
rect 764 156 766 159
rect 665 153 671 155
rect 659 147 665 149
rect 659 145 661 147
rect 663 145 665 147
rect 659 143 665 145
rect 659 140 661 143
rect 669 140 671 153
rect 679 154 685 156
rect 679 152 681 154
rect 683 152 685 154
rect 679 150 685 152
rect 689 154 711 156
rect 689 152 700 154
rect 702 152 707 154
rect 709 152 711 154
rect 689 150 711 152
rect 715 154 721 156
rect 715 152 717 154
rect 719 152 721 154
rect 715 150 721 152
rect 725 154 731 156
rect 725 152 727 154
rect 729 152 731 154
rect 725 150 731 152
rect 754 154 760 156
rect 754 152 756 154
rect 758 152 760 154
rect 764 153 768 156
rect 754 150 760 152
rect 679 147 681 150
rect 689 147 691 150
rect 709 147 711 150
rect 716 147 718 150
rect 619 132 621 136
rect 629 132 631 136
rect 639 132 641 136
rect 580 123 582 127
rect 587 123 589 127
rect 598 123 600 127
rect 659 123 661 127
rect 669 125 671 130
rect 679 128 681 133
rect 689 128 691 133
rect 727 141 729 150
rect 754 142 756 150
rect 766 139 768 153
rect 774 148 776 159
rect 773 146 779 148
rect 773 144 775 146
rect 777 144 779 146
rect 773 142 779 144
rect 773 139 775 142
rect 754 132 756 136
rect 709 123 711 127
rect 716 123 718 127
rect 727 123 729 127
rect 766 125 768 130
rect 773 125 775 130
rect 125 93 127 97
rect 91 84 97 86
rect 91 82 93 84
rect 95 82 97 84
rect 81 77 83 82
rect 91 80 97 82
rect 91 75 93 80
rect 101 75 103 80
rect 148 90 150 95
rect 155 90 157 95
rect 173 93 175 97
rect 183 93 185 97
rect 193 93 195 97
rect 138 81 140 86
rect 81 62 83 65
rect 91 62 93 65
rect 81 60 87 62
rect 81 58 83 60
rect 85 58 87 60
rect 91 59 95 62
rect 81 56 87 58
rect 81 48 83 56
rect 93 45 95 59
rect 101 54 103 65
rect 125 55 127 68
rect 138 65 140 68
rect 227 93 229 97
rect 234 93 236 97
rect 254 93 256 97
rect 214 84 216 88
rect 131 63 140 65
rect 131 61 133 63
rect 135 61 137 63
rect 148 62 150 65
rect 155 62 157 65
rect 173 62 175 65
rect 183 62 185 65
rect 193 62 195 65
rect 214 63 216 72
rect 227 70 229 75
rect 224 68 230 70
rect 224 66 226 68
rect 228 66 230 68
rect 224 64 230 66
rect 131 59 137 61
rect 100 52 106 54
rect 100 50 102 52
rect 104 50 106 52
rect 100 48 106 50
rect 125 53 131 55
rect 125 51 127 53
rect 129 51 131 53
rect 125 49 131 51
rect 100 45 102 48
rect 125 46 127 49
rect 135 46 137 59
rect 145 60 151 62
rect 145 58 147 60
rect 149 58 151 60
rect 145 56 151 58
rect 155 60 177 62
rect 155 58 166 60
rect 168 58 173 60
rect 175 58 177 60
rect 155 56 177 58
rect 181 60 187 62
rect 181 58 183 60
rect 185 58 187 60
rect 181 56 187 58
rect 191 60 197 62
rect 191 58 193 60
rect 195 58 197 60
rect 191 56 197 58
rect 214 61 220 63
rect 214 59 216 61
rect 218 59 220 61
rect 214 57 220 59
rect 145 53 147 56
rect 155 53 157 56
rect 175 53 177 56
rect 182 53 184 56
rect 81 38 83 42
rect 93 31 95 36
rect 100 31 102 36
rect 125 29 127 33
rect 135 31 137 36
rect 145 34 147 39
rect 155 34 157 39
rect 193 47 195 56
rect 214 48 216 57
rect 224 48 226 64
rect 234 62 236 75
rect 277 90 279 95
rect 284 90 286 95
rect 302 93 304 97
rect 312 93 314 97
rect 322 93 324 97
rect 267 81 269 86
rect 234 60 240 62
rect 234 58 236 60
rect 238 58 240 60
rect 234 56 240 58
rect 234 48 236 56
rect 254 55 256 68
rect 267 65 269 68
rect 391 93 393 97
rect 358 84 364 86
rect 358 82 360 84
rect 362 82 364 84
rect 348 77 350 82
rect 358 80 364 82
rect 358 75 360 80
rect 368 75 370 80
rect 414 90 416 95
rect 421 90 423 95
rect 439 93 441 97
rect 449 93 451 97
rect 459 93 461 97
rect 404 81 406 86
rect 260 63 269 65
rect 260 61 262 63
rect 264 61 266 63
rect 277 62 279 65
rect 284 62 286 65
rect 302 62 304 65
rect 312 62 314 65
rect 322 62 324 65
rect 348 62 350 65
rect 358 62 360 65
rect 260 59 266 61
rect 254 53 260 55
rect 254 51 256 53
rect 258 51 260 53
rect 254 49 260 51
rect 254 46 256 49
rect 264 46 266 59
rect 274 60 280 62
rect 274 58 276 60
rect 278 58 280 60
rect 274 56 280 58
rect 284 60 306 62
rect 284 58 295 60
rect 297 58 302 60
rect 304 58 306 60
rect 284 56 306 58
rect 310 60 316 62
rect 310 58 312 60
rect 314 58 316 60
rect 310 56 316 58
rect 320 60 326 62
rect 320 58 322 60
rect 324 58 326 60
rect 320 56 326 58
rect 348 60 354 62
rect 348 58 350 60
rect 352 58 354 60
rect 358 59 362 62
rect 348 56 354 58
rect 274 53 276 56
rect 284 53 286 56
rect 304 53 306 56
rect 311 53 313 56
rect 214 38 216 42
rect 224 38 226 42
rect 234 38 236 42
rect 175 29 177 33
rect 182 29 184 33
rect 193 29 195 33
rect 254 29 256 33
rect 264 31 266 36
rect 274 34 276 39
rect 284 34 286 39
rect 322 47 324 56
rect 348 48 350 56
rect 360 45 362 59
rect 368 54 370 65
rect 391 55 393 68
rect 404 65 406 68
rect 493 93 495 97
rect 500 93 502 97
rect 520 93 522 97
rect 480 84 482 88
rect 397 63 406 65
rect 397 61 399 63
rect 401 61 403 63
rect 414 62 416 65
rect 421 62 423 65
rect 439 62 441 65
rect 449 62 451 65
rect 459 62 461 65
rect 480 63 482 72
rect 493 70 495 75
rect 490 68 496 70
rect 490 66 492 68
rect 494 66 496 68
rect 490 64 496 66
rect 397 59 403 61
rect 367 52 373 54
rect 367 50 369 52
rect 371 50 373 52
rect 367 48 373 50
rect 391 53 397 55
rect 391 51 393 53
rect 395 51 397 53
rect 391 49 397 51
rect 367 45 369 48
rect 391 46 393 49
rect 401 46 403 59
rect 411 60 417 62
rect 411 58 413 60
rect 415 58 417 60
rect 411 56 417 58
rect 421 60 443 62
rect 421 58 432 60
rect 434 58 439 60
rect 441 58 443 60
rect 421 56 443 58
rect 447 60 453 62
rect 447 58 449 60
rect 451 58 453 60
rect 447 56 453 58
rect 457 60 463 62
rect 457 58 459 60
rect 461 58 463 60
rect 457 56 463 58
rect 480 61 486 63
rect 480 59 482 61
rect 484 59 486 61
rect 480 57 486 59
rect 411 53 413 56
rect 421 53 423 56
rect 441 53 443 56
rect 448 53 450 56
rect 348 38 350 42
rect 304 29 306 33
rect 311 29 313 33
rect 322 29 324 33
rect 360 31 362 36
rect 367 31 369 36
rect 391 29 393 33
rect 401 31 403 36
rect 411 34 413 39
rect 421 34 423 39
rect 459 47 461 56
rect 480 48 482 57
rect 490 48 492 64
rect 500 62 502 75
rect 543 90 545 95
rect 550 90 552 95
rect 568 93 570 97
rect 578 93 580 97
rect 588 93 590 97
rect 533 81 535 86
rect 500 60 506 62
rect 500 58 502 60
rect 504 58 506 60
rect 500 56 506 58
rect 500 48 502 56
rect 520 55 522 68
rect 533 65 535 68
rect 657 93 659 97
rect 625 84 631 86
rect 625 82 627 84
rect 629 82 631 84
rect 615 77 617 82
rect 625 80 631 82
rect 625 75 627 80
rect 635 75 637 80
rect 680 90 682 95
rect 687 90 689 95
rect 705 93 707 97
rect 715 93 717 97
rect 725 93 727 97
rect 670 81 672 86
rect 526 63 535 65
rect 526 61 528 63
rect 530 61 532 63
rect 543 62 545 65
rect 550 62 552 65
rect 568 62 570 65
rect 578 62 580 65
rect 588 62 590 65
rect 615 62 617 65
rect 625 62 627 65
rect 526 59 532 61
rect 520 53 526 55
rect 520 51 522 53
rect 524 51 526 53
rect 520 49 526 51
rect 520 46 522 49
rect 530 46 532 59
rect 540 60 546 62
rect 540 58 542 60
rect 544 58 546 60
rect 540 56 546 58
rect 550 60 572 62
rect 550 58 561 60
rect 563 58 568 60
rect 570 58 572 60
rect 550 56 572 58
rect 576 60 582 62
rect 576 58 578 60
rect 580 58 582 60
rect 576 56 582 58
rect 586 60 592 62
rect 586 58 588 60
rect 590 58 592 60
rect 586 56 592 58
rect 615 60 621 62
rect 615 58 617 60
rect 619 58 621 60
rect 625 59 629 62
rect 615 56 621 58
rect 540 53 542 56
rect 550 53 552 56
rect 570 53 572 56
rect 577 53 579 56
rect 480 38 482 42
rect 490 38 492 42
rect 500 38 502 42
rect 441 29 443 33
rect 448 29 450 33
rect 459 29 461 33
rect 520 29 522 33
rect 530 31 532 36
rect 540 34 542 39
rect 550 34 552 39
rect 588 47 590 56
rect 615 48 617 56
rect 627 45 629 59
rect 635 54 637 65
rect 657 55 659 68
rect 670 65 672 68
rect 759 93 761 97
rect 766 93 768 97
rect 786 93 788 97
rect 746 84 748 88
rect 663 63 672 65
rect 663 61 665 63
rect 667 61 669 63
rect 680 62 682 65
rect 687 62 689 65
rect 705 62 707 65
rect 715 62 717 65
rect 725 62 727 65
rect 746 63 748 72
rect 759 70 761 75
rect 756 68 762 70
rect 756 66 758 68
rect 760 66 762 68
rect 756 64 762 66
rect 663 59 669 61
rect 634 52 640 54
rect 634 50 636 52
rect 638 50 640 52
rect 634 48 640 50
rect 657 53 663 55
rect 657 51 659 53
rect 661 51 663 53
rect 657 49 663 51
rect 634 45 636 48
rect 657 46 659 49
rect 667 46 669 59
rect 677 60 683 62
rect 677 58 679 60
rect 681 58 683 60
rect 677 56 683 58
rect 687 60 709 62
rect 687 58 698 60
rect 700 58 705 60
rect 707 58 709 60
rect 687 56 709 58
rect 713 60 719 62
rect 713 58 715 60
rect 717 58 719 60
rect 713 56 719 58
rect 723 60 729 62
rect 723 58 725 60
rect 727 58 729 60
rect 723 56 729 58
rect 746 61 752 63
rect 746 59 748 61
rect 750 59 752 61
rect 746 57 752 59
rect 677 53 679 56
rect 687 53 689 56
rect 707 53 709 56
rect 714 53 716 56
rect 615 38 617 42
rect 570 29 572 33
rect 577 29 579 33
rect 588 29 590 33
rect 627 31 629 36
rect 634 31 636 36
rect 657 29 659 33
rect 667 31 669 36
rect 677 34 679 39
rect 687 34 689 39
rect 725 47 727 56
rect 746 48 748 57
rect 756 48 758 64
rect 766 62 768 75
rect 809 90 811 95
rect 816 90 818 95
rect 834 93 836 97
rect 844 93 846 97
rect 854 93 856 97
rect 799 81 801 86
rect 766 60 772 62
rect 766 58 768 60
rect 770 58 772 60
rect 766 56 772 58
rect 766 48 768 56
rect 786 55 788 68
rect 799 65 801 68
rect 890 84 896 86
rect 890 82 892 84
rect 894 82 896 84
rect 880 77 882 82
rect 890 80 896 82
rect 890 75 892 80
rect 900 75 902 80
rect 792 63 801 65
rect 792 61 794 63
rect 796 61 798 63
rect 809 62 811 65
rect 816 62 818 65
rect 834 62 836 65
rect 844 62 846 65
rect 854 62 856 65
rect 880 62 882 65
rect 890 62 892 65
rect 792 59 798 61
rect 786 53 792 55
rect 786 51 788 53
rect 790 51 792 53
rect 786 49 792 51
rect 786 46 788 49
rect 796 46 798 59
rect 806 60 812 62
rect 806 58 808 60
rect 810 58 812 60
rect 806 56 812 58
rect 816 60 838 62
rect 816 58 827 60
rect 829 58 834 60
rect 836 58 838 60
rect 816 56 838 58
rect 842 60 848 62
rect 842 58 844 60
rect 846 58 848 60
rect 842 56 848 58
rect 852 60 858 62
rect 852 58 854 60
rect 856 58 858 60
rect 852 56 858 58
rect 880 60 886 62
rect 880 58 882 60
rect 884 58 886 60
rect 890 59 894 62
rect 880 56 886 58
rect 806 53 808 56
rect 816 53 818 56
rect 836 53 838 56
rect 843 53 845 56
rect 746 38 748 42
rect 756 38 758 42
rect 766 38 768 42
rect 707 29 709 33
rect 714 29 716 33
rect 725 29 727 33
rect 786 29 788 33
rect 796 31 798 36
rect 806 34 808 39
rect 816 34 818 39
rect 854 47 856 56
rect 880 48 882 56
rect 892 45 894 59
rect 900 54 902 65
rect 899 52 905 54
rect 899 50 901 52
rect 903 50 905 52
rect 899 48 905 50
rect 899 45 901 48
rect 880 38 882 42
rect 836 29 838 33
rect 843 29 845 33
rect 854 29 856 33
rect 892 31 894 36
rect 899 31 901 36
<< ndif >>
rect 97 328 102 335
rect 75 326 82 328
rect 75 324 77 326
rect 79 324 82 326
rect 75 322 82 324
rect 77 315 82 322
rect 84 322 92 328
rect 84 320 87 322
rect 89 320 92 322
rect 84 318 92 320
rect 94 325 102 328
rect 94 323 97 325
rect 99 323 102 325
rect 94 321 102 323
rect 104 333 112 335
rect 104 331 107 333
rect 109 331 112 333
rect 104 321 112 331
rect 114 333 121 335
rect 114 331 117 333
rect 119 331 121 333
rect 114 326 121 331
rect 127 328 132 335
rect 114 324 117 326
rect 119 324 121 326
rect 114 321 121 324
rect 125 326 132 328
rect 125 324 127 326
rect 129 324 132 326
rect 125 322 132 324
rect 94 318 99 321
rect 84 315 89 318
rect 127 315 132 322
rect 134 315 139 335
rect 141 329 148 335
rect 141 319 150 329
rect 141 317 144 319
rect 146 317 150 319
rect 141 315 150 317
rect 152 326 164 329
rect 197 328 202 335
rect 152 324 155 326
rect 157 324 164 326
rect 152 315 164 324
rect 175 326 182 328
rect 175 324 177 326
rect 179 324 182 326
rect 175 322 182 324
rect 177 315 182 322
rect 184 322 192 328
rect 184 320 187 322
rect 189 320 192 322
rect 184 318 192 320
rect 194 325 202 328
rect 194 323 197 325
rect 199 323 202 325
rect 194 321 202 323
rect 204 333 212 335
rect 204 331 207 333
rect 209 331 212 333
rect 204 321 212 331
rect 214 333 221 335
rect 214 331 217 333
rect 219 331 221 333
rect 214 326 221 331
rect 227 328 232 335
rect 214 324 217 326
rect 219 324 221 326
rect 214 321 221 324
rect 225 326 232 328
rect 225 324 227 326
rect 229 324 232 326
rect 225 322 232 324
rect 194 318 199 321
rect 184 315 189 318
rect 227 315 232 322
rect 234 315 239 335
rect 241 329 248 335
rect 241 319 250 329
rect 241 317 244 319
rect 246 317 250 319
rect 241 315 250 317
rect 252 326 259 329
rect 252 324 255 326
rect 257 324 259 326
rect 264 328 271 330
rect 264 326 266 328
rect 268 326 271 328
rect 264 324 271 326
rect 273 328 281 330
rect 273 326 276 328
rect 278 326 281 328
rect 273 324 281 326
rect 283 328 291 330
rect 283 326 286 328
rect 288 326 291 328
rect 283 324 291 326
rect 293 328 300 330
rect 326 328 331 335
rect 293 326 296 328
rect 298 326 300 328
rect 293 324 300 326
rect 304 326 311 328
rect 304 324 306 326
rect 308 324 311 326
rect 252 322 259 324
rect 252 315 257 322
rect 304 322 311 324
rect 306 315 311 322
rect 313 322 321 328
rect 313 320 316 322
rect 318 320 321 322
rect 313 318 321 320
rect 323 325 331 328
rect 323 323 326 325
rect 328 323 331 325
rect 323 321 331 323
rect 333 333 341 335
rect 333 331 336 333
rect 338 331 341 333
rect 333 321 341 331
rect 343 333 350 335
rect 343 331 346 333
rect 348 331 350 333
rect 343 326 350 331
rect 356 328 361 335
rect 343 324 346 326
rect 348 324 350 326
rect 343 321 350 324
rect 354 326 361 328
rect 354 324 356 326
rect 358 324 361 326
rect 354 322 361 324
rect 323 318 328 321
rect 313 315 318 318
rect 356 315 361 322
rect 363 315 368 335
rect 370 329 377 335
rect 370 319 379 329
rect 370 317 373 319
rect 375 317 379 319
rect 370 315 379 317
rect 381 326 388 329
rect 421 328 426 335
rect 381 324 384 326
rect 386 324 388 326
rect 381 322 388 324
rect 399 326 406 328
rect 399 324 401 326
rect 403 324 406 326
rect 399 322 406 324
rect 381 315 386 322
rect 401 315 406 322
rect 408 322 416 328
rect 408 320 411 322
rect 413 320 416 322
rect 408 318 416 320
rect 418 325 426 328
rect 418 323 421 325
rect 423 323 426 325
rect 418 321 426 323
rect 428 333 436 335
rect 428 331 431 333
rect 433 331 436 333
rect 428 321 436 331
rect 438 333 445 335
rect 438 331 441 333
rect 443 331 445 333
rect 438 326 445 331
rect 451 328 456 335
rect 438 324 441 326
rect 443 324 445 326
rect 438 321 445 324
rect 449 326 456 328
rect 449 324 451 326
rect 453 324 456 326
rect 449 322 456 324
rect 418 318 423 321
rect 408 315 413 318
rect 451 315 456 322
rect 458 315 463 335
rect 465 329 472 335
rect 465 319 474 329
rect 465 317 468 319
rect 470 317 474 319
rect 465 315 474 317
rect 476 326 483 329
rect 476 324 479 326
rect 481 324 483 326
rect 488 328 495 330
rect 488 326 490 328
rect 492 326 495 328
rect 488 324 495 326
rect 497 328 505 330
rect 497 326 500 328
rect 502 326 505 328
rect 497 324 505 326
rect 507 328 515 330
rect 507 326 510 328
rect 512 326 515 328
rect 507 324 515 326
rect 517 328 524 330
rect 550 328 555 335
rect 517 326 520 328
rect 522 326 524 328
rect 517 324 524 326
rect 528 326 535 328
rect 528 324 530 326
rect 532 324 535 326
rect 476 322 483 324
rect 476 315 481 322
rect 528 322 535 324
rect 530 315 535 322
rect 537 322 545 328
rect 537 320 540 322
rect 542 320 545 322
rect 537 318 545 320
rect 547 325 555 328
rect 547 323 550 325
rect 552 323 555 325
rect 547 321 555 323
rect 557 333 565 335
rect 557 331 560 333
rect 562 331 565 333
rect 557 321 565 331
rect 567 333 574 335
rect 567 331 570 333
rect 572 331 574 333
rect 567 326 574 331
rect 580 328 585 335
rect 567 324 570 326
rect 572 324 574 326
rect 567 321 574 324
rect 578 326 585 328
rect 578 324 580 326
rect 582 324 585 326
rect 578 322 585 324
rect 547 318 552 321
rect 537 315 542 318
rect 580 315 585 322
rect 587 315 592 335
rect 594 329 601 335
rect 594 319 603 329
rect 594 317 597 319
rect 599 317 603 319
rect 594 315 603 317
rect 605 326 612 329
rect 646 328 651 335
rect 605 324 608 326
rect 610 324 612 326
rect 605 322 612 324
rect 624 326 631 328
rect 624 324 626 326
rect 628 324 631 326
rect 624 322 631 324
rect 605 315 610 322
rect 626 315 631 322
rect 633 322 641 328
rect 633 320 636 322
rect 638 320 641 322
rect 633 318 641 320
rect 643 325 651 328
rect 643 323 646 325
rect 648 323 651 325
rect 643 321 651 323
rect 653 333 661 335
rect 653 331 656 333
rect 658 331 661 333
rect 653 321 661 331
rect 663 333 670 335
rect 663 331 666 333
rect 668 331 670 333
rect 663 326 670 331
rect 676 328 681 335
rect 663 324 666 326
rect 668 324 670 326
rect 663 321 670 324
rect 674 326 681 328
rect 674 324 676 326
rect 678 324 681 326
rect 674 322 681 324
rect 643 318 648 321
rect 633 315 638 318
rect 676 315 681 322
rect 683 315 688 335
rect 690 329 697 335
rect 690 319 699 329
rect 690 317 693 319
rect 695 317 699 319
rect 690 315 699 317
rect 701 326 708 329
rect 701 324 704 326
rect 706 324 708 326
rect 723 328 730 330
rect 723 326 725 328
rect 727 326 730 328
rect 723 324 730 326
rect 732 327 740 330
rect 772 328 779 330
rect 732 324 742 327
rect 701 322 708 324
rect 701 315 706 322
rect 734 318 742 324
rect 744 318 749 327
rect 751 325 758 327
rect 751 323 754 325
rect 756 323 758 325
rect 772 326 774 328
rect 776 326 779 328
rect 772 324 779 326
rect 781 327 789 330
rect 822 328 829 330
rect 781 324 791 327
rect 751 321 758 323
rect 751 318 756 321
rect 783 318 791 324
rect 793 318 798 327
rect 800 325 807 327
rect 800 323 803 325
rect 805 323 807 325
rect 822 326 824 328
rect 826 326 829 328
rect 822 324 829 326
rect 831 327 839 330
rect 831 324 841 327
rect 800 321 807 323
rect 800 318 805 321
rect 833 318 841 324
rect 843 318 848 327
rect 850 325 857 327
rect 850 323 853 325
rect 855 323 857 325
rect 850 321 857 323
rect 850 318 855 321
rect 734 316 740 318
rect 734 314 736 316
rect 738 314 740 316
rect 734 312 740 314
rect 783 316 789 318
rect 783 314 785 316
rect 787 314 789 316
rect 783 312 789 314
rect 833 316 839 318
rect 833 314 835 316
rect 837 314 839 316
rect 833 312 839 314
rect 75 234 82 236
rect 75 232 77 234
rect 79 232 82 234
rect 75 230 82 232
rect 84 233 92 236
rect 125 234 132 236
rect 84 230 94 233
rect 86 224 94 230
rect 96 224 101 233
rect 103 231 110 233
rect 103 229 106 231
rect 108 229 110 231
rect 125 232 127 234
rect 129 232 132 234
rect 125 230 132 232
rect 134 233 142 236
rect 196 235 203 237
rect 196 233 198 235
rect 200 233 203 235
rect 134 230 144 233
rect 103 227 110 229
rect 103 224 108 227
rect 136 224 144 230
rect 146 224 151 233
rect 153 231 160 233
rect 196 231 203 233
rect 205 234 213 237
rect 237 235 244 237
rect 205 231 215 234
rect 153 229 156 231
rect 158 229 160 231
rect 153 227 160 229
rect 153 224 158 227
rect 207 225 215 231
rect 217 225 222 234
rect 224 232 231 234
rect 224 230 227 232
rect 229 230 231 232
rect 237 233 239 235
rect 241 233 244 235
rect 237 231 244 233
rect 246 234 254 237
rect 325 234 332 236
rect 246 231 256 234
rect 224 228 231 230
rect 224 225 229 228
rect 248 225 256 231
rect 258 225 263 234
rect 265 232 272 234
rect 265 230 268 232
rect 270 230 272 232
rect 325 232 327 234
rect 329 232 332 234
rect 325 230 332 232
rect 334 233 342 236
rect 375 234 382 236
rect 334 230 344 233
rect 265 228 272 230
rect 265 225 270 228
rect 86 222 92 224
rect 86 220 88 222
rect 90 220 92 222
rect 86 218 92 220
rect 136 222 142 224
rect 136 220 138 222
rect 140 220 142 222
rect 136 218 142 220
rect 207 223 213 225
rect 207 221 209 223
rect 211 221 213 223
rect 207 219 213 221
rect 248 223 254 225
rect 248 221 250 223
rect 252 221 254 223
rect 248 219 254 221
rect 336 224 344 230
rect 346 224 351 233
rect 353 231 360 233
rect 353 229 356 231
rect 358 229 360 231
rect 375 232 377 234
rect 379 232 382 234
rect 375 230 382 232
rect 384 233 392 236
rect 419 234 426 236
rect 384 230 394 233
rect 353 227 360 229
rect 353 224 358 227
rect 386 224 394 230
rect 396 224 401 233
rect 403 231 410 233
rect 403 229 406 231
rect 408 229 410 231
rect 419 232 421 234
rect 423 232 426 234
rect 419 230 426 232
rect 428 233 436 236
rect 475 234 482 236
rect 428 230 438 233
rect 403 227 410 229
rect 403 224 408 227
rect 430 224 438 230
rect 440 224 445 233
rect 447 231 454 233
rect 447 229 450 231
rect 452 229 454 231
rect 475 232 477 234
rect 479 232 482 234
rect 475 230 482 232
rect 484 233 492 236
rect 525 234 532 236
rect 484 230 494 233
rect 447 227 454 229
rect 447 224 452 227
rect 486 224 494 230
rect 496 224 501 233
rect 503 231 510 233
rect 503 229 506 231
rect 508 229 510 231
rect 525 232 527 234
rect 529 232 532 234
rect 525 230 532 232
rect 534 233 542 236
rect 575 234 582 236
rect 534 230 544 233
rect 503 227 510 229
rect 503 224 508 227
rect 536 224 544 230
rect 546 224 551 233
rect 553 231 560 233
rect 553 229 556 231
rect 558 229 560 231
rect 575 232 577 234
rect 579 232 582 234
rect 575 230 582 232
rect 584 233 592 236
rect 625 234 632 236
rect 584 230 594 233
rect 553 227 560 229
rect 553 224 558 227
rect 586 224 594 230
rect 596 224 601 233
rect 603 231 610 233
rect 603 229 606 231
rect 608 229 610 231
rect 625 232 627 234
rect 629 232 632 234
rect 625 230 632 232
rect 634 233 642 236
rect 691 234 696 241
rect 634 230 644 233
rect 603 227 610 229
rect 603 224 608 227
rect 636 224 644 230
rect 646 224 651 233
rect 653 231 660 233
rect 653 229 656 231
rect 658 229 660 231
rect 653 227 660 229
rect 669 232 676 234
rect 669 230 671 232
rect 673 230 676 232
rect 669 228 676 230
rect 653 224 658 227
rect 336 222 342 224
rect 336 220 338 222
rect 340 220 342 222
rect 336 218 342 220
rect 386 222 392 224
rect 386 220 388 222
rect 390 220 392 222
rect 386 218 392 220
rect 430 222 436 224
rect 430 220 432 222
rect 434 220 436 222
rect 430 218 436 220
rect 486 222 492 224
rect 486 220 488 222
rect 490 220 492 222
rect 486 218 492 220
rect 536 222 542 224
rect 536 220 538 222
rect 540 220 542 222
rect 536 218 542 220
rect 586 222 592 224
rect 586 220 588 222
rect 590 220 592 222
rect 586 218 592 220
rect 636 222 642 224
rect 636 220 638 222
rect 640 220 642 222
rect 636 218 642 220
rect 671 221 676 228
rect 678 228 686 234
rect 678 226 681 228
rect 683 226 686 228
rect 678 224 686 226
rect 688 231 696 234
rect 688 229 691 231
rect 693 229 696 231
rect 688 227 696 229
rect 698 239 706 241
rect 698 237 701 239
rect 703 237 706 239
rect 698 227 706 237
rect 708 239 715 241
rect 708 237 711 239
rect 713 237 715 239
rect 708 232 715 237
rect 721 234 726 241
rect 708 230 711 232
rect 713 230 715 232
rect 708 227 715 230
rect 719 232 726 234
rect 719 230 721 232
rect 723 230 726 232
rect 719 228 726 230
rect 688 224 693 227
rect 678 221 683 224
rect 721 221 726 228
rect 728 221 733 241
rect 735 235 742 241
rect 735 225 744 235
rect 735 223 738 225
rect 740 223 744 225
rect 735 221 744 223
rect 746 232 753 235
rect 791 234 796 241
rect 746 230 749 232
rect 751 230 753 232
rect 746 228 753 230
rect 769 232 776 234
rect 769 230 771 232
rect 773 230 776 232
rect 769 228 776 230
rect 746 221 751 228
rect 771 221 776 228
rect 778 228 786 234
rect 778 226 781 228
rect 783 226 786 228
rect 778 224 786 226
rect 788 231 796 234
rect 788 229 791 231
rect 793 229 796 231
rect 788 227 796 229
rect 798 239 806 241
rect 798 237 801 239
rect 803 237 806 239
rect 798 227 806 237
rect 808 239 815 241
rect 808 237 811 239
rect 813 237 815 239
rect 808 232 815 237
rect 821 234 826 241
rect 808 230 811 232
rect 813 230 815 232
rect 808 227 815 230
rect 819 232 826 234
rect 819 230 821 232
rect 823 230 826 232
rect 819 228 826 230
rect 788 224 793 227
rect 778 221 783 224
rect 821 221 826 228
rect 828 221 833 241
rect 835 235 842 241
rect 835 225 844 235
rect 835 223 838 225
rect 840 223 844 225
rect 835 221 844 223
rect 846 232 853 235
rect 846 230 849 232
rect 851 230 853 232
rect 846 228 853 230
rect 846 221 851 228
rect 97 140 102 147
rect 75 138 82 140
rect 75 136 77 138
rect 79 136 82 138
rect 75 134 82 136
rect 77 127 82 134
rect 84 134 92 140
rect 84 132 87 134
rect 89 132 92 134
rect 84 130 92 132
rect 94 137 102 140
rect 94 135 97 137
rect 99 135 102 137
rect 94 133 102 135
rect 104 145 112 147
rect 104 143 107 145
rect 109 143 112 145
rect 104 133 112 143
rect 114 145 121 147
rect 114 143 117 145
rect 119 143 121 145
rect 114 138 121 143
rect 127 140 132 147
rect 114 136 117 138
rect 119 136 121 138
rect 114 133 121 136
rect 125 138 132 140
rect 125 136 127 138
rect 129 136 132 138
rect 125 134 132 136
rect 94 130 99 133
rect 84 127 89 130
rect 127 127 132 134
rect 134 127 139 147
rect 141 141 148 147
rect 141 131 150 141
rect 141 129 144 131
rect 146 129 150 131
rect 141 127 150 129
rect 152 138 159 141
rect 152 136 155 138
rect 157 136 159 138
rect 164 140 171 142
rect 164 138 166 140
rect 168 138 171 140
rect 164 136 171 138
rect 173 140 181 142
rect 173 138 176 140
rect 178 138 181 140
rect 173 136 181 138
rect 183 140 191 142
rect 183 138 186 140
rect 188 138 191 140
rect 183 136 191 138
rect 193 140 200 142
rect 226 140 231 147
rect 193 138 196 140
rect 198 138 200 140
rect 193 136 200 138
rect 204 138 211 140
rect 204 136 206 138
rect 208 136 211 138
rect 152 134 159 136
rect 152 127 157 134
rect 204 134 211 136
rect 206 127 211 134
rect 213 134 221 140
rect 213 132 216 134
rect 218 132 221 134
rect 213 130 221 132
rect 223 137 231 140
rect 223 135 226 137
rect 228 135 231 137
rect 223 133 231 135
rect 233 145 241 147
rect 233 143 236 145
rect 238 143 241 145
rect 233 133 241 143
rect 243 145 250 147
rect 243 143 246 145
rect 248 143 250 145
rect 243 138 250 143
rect 256 140 261 147
rect 243 136 246 138
rect 248 136 250 138
rect 243 133 250 136
rect 254 138 261 140
rect 254 136 256 138
rect 258 136 261 138
rect 254 134 261 136
rect 223 130 228 133
rect 213 127 218 130
rect 256 127 261 134
rect 263 127 268 147
rect 270 141 277 147
rect 270 131 279 141
rect 270 129 273 131
rect 275 129 279 131
rect 270 127 279 129
rect 281 138 288 141
rect 281 136 284 138
rect 286 136 288 138
rect 281 134 288 136
rect 298 140 303 146
rect 321 140 326 147
rect 281 127 286 134
rect 298 127 306 140
rect 308 134 316 140
rect 308 132 311 134
rect 313 132 316 134
rect 308 130 316 132
rect 318 137 326 140
rect 318 135 321 137
rect 323 135 326 137
rect 318 133 326 135
rect 328 145 336 147
rect 328 143 331 145
rect 333 143 336 145
rect 328 133 336 143
rect 338 145 345 147
rect 338 143 341 145
rect 343 143 345 145
rect 338 138 345 143
rect 351 140 356 147
rect 338 136 341 138
rect 343 136 345 138
rect 338 133 345 136
rect 349 138 356 140
rect 349 136 351 138
rect 353 136 356 138
rect 349 134 356 136
rect 318 130 323 133
rect 308 127 313 130
rect 298 120 304 127
rect 351 127 356 134
rect 358 127 363 147
rect 365 141 372 147
rect 365 131 374 141
rect 365 129 368 131
rect 370 129 374 131
rect 365 127 374 129
rect 376 138 383 141
rect 376 136 379 138
rect 381 136 383 138
rect 388 140 395 142
rect 388 138 390 140
rect 392 138 395 140
rect 388 136 395 138
rect 397 140 405 142
rect 397 138 400 140
rect 402 138 405 140
rect 397 136 405 138
rect 407 140 415 142
rect 407 138 410 140
rect 412 138 415 140
rect 407 136 415 138
rect 417 140 424 142
rect 450 140 455 147
rect 417 138 420 140
rect 422 138 424 140
rect 417 136 424 138
rect 428 138 435 140
rect 428 136 430 138
rect 432 136 435 138
rect 376 134 383 136
rect 376 127 381 134
rect 428 134 435 136
rect 430 127 435 134
rect 437 134 445 140
rect 437 132 440 134
rect 442 132 445 134
rect 437 130 445 132
rect 447 137 455 140
rect 447 135 450 137
rect 452 135 455 137
rect 447 133 455 135
rect 457 145 465 147
rect 457 143 460 145
rect 462 143 465 145
rect 457 133 465 143
rect 467 145 474 147
rect 467 143 470 145
rect 472 143 474 145
rect 467 138 474 143
rect 480 140 485 147
rect 467 136 470 138
rect 472 136 474 138
rect 467 133 474 136
rect 478 138 485 140
rect 478 136 480 138
rect 482 136 485 138
rect 478 134 485 136
rect 447 130 452 133
rect 437 127 442 130
rect 480 127 485 134
rect 487 127 492 147
rect 494 141 501 147
rect 494 131 503 141
rect 494 129 497 131
rect 499 129 503 131
rect 494 127 503 129
rect 505 138 512 141
rect 545 140 550 147
rect 505 136 508 138
rect 510 136 512 138
rect 505 134 512 136
rect 523 138 530 140
rect 523 136 525 138
rect 527 136 530 138
rect 523 134 530 136
rect 505 127 510 134
rect 525 127 530 134
rect 532 134 540 140
rect 532 132 535 134
rect 537 132 540 134
rect 532 130 540 132
rect 542 137 550 140
rect 542 135 545 137
rect 547 135 550 137
rect 542 133 550 135
rect 552 145 560 147
rect 552 143 555 145
rect 557 143 560 145
rect 552 133 560 143
rect 562 145 569 147
rect 562 143 565 145
rect 567 143 569 145
rect 562 138 569 143
rect 575 140 580 147
rect 562 136 565 138
rect 567 136 569 138
rect 562 133 569 136
rect 573 138 580 140
rect 573 136 575 138
rect 577 136 580 138
rect 573 134 580 136
rect 542 130 547 133
rect 532 127 537 130
rect 575 127 580 134
rect 582 127 587 147
rect 589 141 596 147
rect 589 131 598 141
rect 589 129 592 131
rect 594 129 598 131
rect 589 127 598 129
rect 600 138 607 141
rect 600 136 603 138
rect 605 136 607 138
rect 612 140 619 142
rect 612 138 614 140
rect 616 138 619 140
rect 612 136 619 138
rect 621 140 629 142
rect 621 138 624 140
rect 626 138 629 140
rect 621 136 629 138
rect 631 140 639 142
rect 631 138 634 140
rect 636 138 639 140
rect 631 136 639 138
rect 641 140 648 142
rect 674 140 679 147
rect 641 138 644 140
rect 646 138 648 140
rect 641 136 648 138
rect 652 138 659 140
rect 652 136 654 138
rect 656 136 659 138
rect 600 134 607 136
rect 600 127 605 134
rect 652 134 659 136
rect 654 127 659 134
rect 661 134 669 140
rect 661 132 664 134
rect 666 132 669 134
rect 661 130 669 132
rect 671 137 679 140
rect 671 135 674 137
rect 676 135 679 137
rect 671 133 679 135
rect 681 145 689 147
rect 681 143 684 145
rect 686 143 689 145
rect 681 133 689 143
rect 691 145 698 147
rect 691 143 694 145
rect 696 143 698 145
rect 691 138 698 143
rect 704 140 709 147
rect 691 136 694 138
rect 696 136 698 138
rect 691 133 698 136
rect 702 138 709 140
rect 702 136 704 138
rect 706 136 709 138
rect 702 134 709 136
rect 671 130 676 133
rect 661 127 666 130
rect 704 127 709 134
rect 711 127 716 147
rect 718 141 725 147
rect 718 131 727 141
rect 718 129 721 131
rect 723 129 727 131
rect 718 127 727 129
rect 729 138 736 141
rect 729 136 732 138
rect 734 136 736 138
rect 747 140 754 142
rect 747 138 749 140
rect 751 138 754 140
rect 747 136 754 138
rect 756 139 764 142
rect 756 136 766 139
rect 729 134 736 136
rect 729 127 734 134
rect 758 130 766 136
rect 768 130 773 139
rect 775 137 782 139
rect 775 135 778 137
rect 780 135 782 137
rect 775 133 782 135
rect 775 130 780 133
rect 758 128 764 130
rect 758 126 760 128
rect 762 126 764 128
rect 758 124 764 126
rect 74 46 81 48
rect 74 44 76 46
rect 78 44 81 46
rect 74 42 81 44
rect 83 45 91 48
rect 140 46 145 53
rect 83 42 93 45
rect 85 36 93 42
rect 95 36 100 45
rect 102 43 109 45
rect 102 41 105 43
rect 107 41 109 43
rect 102 39 109 41
rect 118 44 125 46
rect 118 42 120 44
rect 122 42 125 44
rect 118 40 125 42
rect 102 36 107 39
rect 85 34 91 36
rect 85 32 87 34
rect 89 32 91 34
rect 85 30 91 32
rect 120 33 125 40
rect 127 40 135 46
rect 127 38 130 40
rect 132 38 135 40
rect 127 36 135 38
rect 137 43 145 46
rect 137 41 140 43
rect 142 41 145 43
rect 137 39 145 41
rect 147 51 155 53
rect 147 49 150 51
rect 152 49 155 51
rect 147 39 155 49
rect 157 51 164 53
rect 157 49 160 51
rect 162 49 164 51
rect 157 44 164 49
rect 170 46 175 53
rect 157 42 160 44
rect 162 42 164 44
rect 157 39 164 42
rect 168 44 175 46
rect 168 42 170 44
rect 172 42 175 44
rect 168 40 175 42
rect 137 36 142 39
rect 127 33 132 36
rect 170 33 175 40
rect 177 33 182 53
rect 184 47 191 53
rect 184 37 193 47
rect 184 35 187 37
rect 189 35 193 37
rect 184 33 193 35
rect 195 44 202 47
rect 195 42 198 44
rect 200 42 202 44
rect 207 46 214 48
rect 207 44 209 46
rect 211 44 214 46
rect 207 42 214 44
rect 216 46 224 48
rect 216 44 219 46
rect 221 44 224 46
rect 216 42 224 44
rect 226 46 234 48
rect 226 44 229 46
rect 231 44 234 46
rect 226 42 234 44
rect 236 46 243 48
rect 269 46 274 53
rect 236 44 239 46
rect 241 44 243 46
rect 236 42 243 44
rect 247 44 254 46
rect 247 42 249 44
rect 251 42 254 44
rect 195 40 202 42
rect 195 33 200 40
rect 247 40 254 42
rect 249 33 254 40
rect 256 40 264 46
rect 256 38 259 40
rect 261 38 264 40
rect 256 36 264 38
rect 266 43 274 46
rect 266 41 269 43
rect 271 41 274 43
rect 266 39 274 41
rect 276 51 284 53
rect 276 49 279 51
rect 281 49 284 51
rect 276 39 284 49
rect 286 51 293 53
rect 286 49 289 51
rect 291 49 293 51
rect 286 44 293 49
rect 299 46 304 53
rect 286 42 289 44
rect 291 42 293 44
rect 286 39 293 42
rect 297 44 304 46
rect 297 42 299 44
rect 301 42 304 44
rect 297 40 304 42
rect 266 36 271 39
rect 256 33 261 36
rect 299 33 304 40
rect 306 33 311 53
rect 313 47 320 53
rect 313 37 322 47
rect 313 35 316 37
rect 318 35 322 37
rect 313 33 322 35
rect 324 44 331 47
rect 324 42 327 44
rect 329 42 331 44
rect 341 46 348 48
rect 341 44 343 46
rect 345 44 348 46
rect 341 42 348 44
rect 350 45 358 48
rect 406 46 411 53
rect 350 42 360 45
rect 324 40 331 42
rect 324 33 329 40
rect 352 36 360 42
rect 362 36 367 45
rect 369 43 376 45
rect 369 41 372 43
rect 374 41 376 43
rect 369 39 376 41
rect 384 44 391 46
rect 384 42 386 44
rect 388 42 391 44
rect 384 40 391 42
rect 369 36 374 39
rect 352 34 358 36
rect 352 32 354 34
rect 356 32 358 34
rect 352 30 358 32
rect 386 33 391 40
rect 393 40 401 46
rect 393 38 396 40
rect 398 38 401 40
rect 393 36 401 38
rect 403 43 411 46
rect 403 41 406 43
rect 408 41 411 43
rect 403 39 411 41
rect 413 51 421 53
rect 413 49 416 51
rect 418 49 421 51
rect 413 39 421 49
rect 423 51 430 53
rect 423 49 426 51
rect 428 49 430 51
rect 423 44 430 49
rect 436 46 441 53
rect 423 42 426 44
rect 428 42 430 44
rect 423 39 430 42
rect 434 44 441 46
rect 434 42 436 44
rect 438 42 441 44
rect 434 40 441 42
rect 403 36 408 39
rect 393 33 398 36
rect 436 33 441 40
rect 443 33 448 53
rect 450 47 457 53
rect 450 37 459 47
rect 450 35 453 37
rect 455 35 459 37
rect 450 33 459 35
rect 461 44 468 47
rect 461 42 464 44
rect 466 42 468 44
rect 473 46 480 48
rect 473 44 475 46
rect 477 44 480 46
rect 473 42 480 44
rect 482 46 490 48
rect 482 44 485 46
rect 487 44 490 46
rect 482 42 490 44
rect 492 46 500 48
rect 492 44 495 46
rect 497 44 500 46
rect 492 42 500 44
rect 502 46 509 48
rect 535 46 540 53
rect 502 44 505 46
rect 507 44 509 46
rect 502 42 509 44
rect 513 44 520 46
rect 513 42 515 44
rect 517 42 520 44
rect 461 40 468 42
rect 461 33 466 40
rect 513 40 520 42
rect 515 33 520 40
rect 522 40 530 46
rect 522 38 525 40
rect 527 38 530 40
rect 522 36 530 38
rect 532 43 540 46
rect 532 41 535 43
rect 537 41 540 43
rect 532 39 540 41
rect 542 51 550 53
rect 542 49 545 51
rect 547 49 550 51
rect 542 39 550 49
rect 552 51 559 53
rect 552 49 555 51
rect 557 49 559 51
rect 552 44 559 49
rect 565 46 570 53
rect 552 42 555 44
rect 557 42 559 44
rect 552 39 559 42
rect 563 44 570 46
rect 563 42 565 44
rect 567 42 570 44
rect 563 40 570 42
rect 532 36 537 39
rect 522 33 527 36
rect 565 33 570 40
rect 572 33 577 53
rect 579 47 586 53
rect 579 37 588 47
rect 579 35 582 37
rect 584 35 588 37
rect 579 33 588 35
rect 590 44 597 47
rect 590 42 593 44
rect 595 42 597 44
rect 608 46 615 48
rect 608 44 610 46
rect 612 44 615 46
rect 608 42 615 44
rect 617 45 625 48
rect 672 46 677 53
rect 617 42 627 45
rect 590 40 597 42
rect 590 33 595 40
rect 619 36 627 42
rect 629 36 634 45
rect 636 43 643 45
rect 636 41 639 43
rect 641 41 643 43
rect 636 39 643 41
rect 650 44 657 46
rect 650 42 652 44
rect 654 42 657 44
rect 650 40 657 42
rect 636 36 641 39
rect 619 34 625 36
rect 619 32 621 34
rect 623 32 625 34
rect 619 30 625 32
rect 652 33 657 40
rect 659 40 667 46
rect 659 38 662 40
rect 664 38 667 40
rect 659 36 667 38
rect 669 43 677 46
rect 669 41 672 43
rect 674 41 677 43
rect 669 39 677 41
rect 679 51 687 53
rect 679 49 682 51
rect 684 49 687 51
rect 679 39 687 49
rect 689 51 696 53
rect 689 49 692 51
rect 694 49 696 51
rect 689 44 696 49
rect 702 46 707 53
rect 689 42 692 44
rect 694 42 696 44
rect 689 39 696 42
rect 700 44 707 46
rect 700 42 702 44
rect 704 42 707 44
rect 700 40 707 42
rect 669 36 674 39
rect 659 33 664 36
rect 702 33 707 40
rect 709 33 714 53
rect 716 47 723 53
rect 716 37 725 47
rect 716 35 719 37
rect 721 35 725 37
rect 716 33 725 35
rect 727 44 734 47
rect 727 42 730 44
rect 732 42 734 44
rect 739 46 746 48
rect 739 44 741 46
rect 743 44 746 46
rect 739 42 746 44
rect 748 46 756 48
rect 748 44 751 46
rect 753 44 756 46
rect 748 42 756 44
rect 758 46 766 48
rect 758 44 761 46
rect 763 44 766 46
rect 758 42 766 44
rect 768 46 775 48
rect 801 46 806 53
rect 768 44 771 46
rect 773 44 775 46
rect 768 42 775 44
rect 779 44 786 46
rect 779 42 781 44
rect 783 42 786 44
rect 727 40 734 42
rect 727 33 732 40
rect 779 40 786 42
rect 781 33 786 40
rect 788 40 796 46
rect 788 38 791 40
rect 793 38 796 40
rect 788 36 796 38
rect 798 43 806 46
rect 798 41 801 43
rect 803 41 806 43
rect 798 39 806 41
rect 808 51 816 53
rect 808 49 811 51
rect 813 49 816 51
rect 808 39 816 49
rect 818 51 825 53
rect 818 49 821 51
rect 823 49 825 51
rect 818 44 825 49
rect 831 46 836 53
rect 818 42 821 44
rect 823 42 825 44
rect 818 39 825 42
rect 829 44 836 46
rect 829 42 831 44
rect 833 42 836 44
rect 829 40 836 42
rect 798 36 803 39
rect 788 33 793 36
rect 831 33 836 40
rect 838 33 843 53
rect 845 47 852 53
rect 845 37 854 47
rect 845 35 848 37
rect 850 35 854 37
rect 845 33 854 35
rect 856 44 863 47
rect 856 42 859 44
rect 861 42 863 44
rect 873 46 880 48
rect 873 44 875 46
rect 877 44 880 46
rect 873 42 880 44
rect 882 45 890 48
rect 882 42 892 45
rect 856 40 863 42
rect 856 33 861 40
rect 884 36 892 42
rect 894 36 899 45
rect 901 43 908 45
rect 901 41 904 43
rect 906 41 908 43
rect 901 39 908 41
rect 901 36 906 39
rect 884 34 890 36
rect 884 32 886 34
rect 888 32 890 34
rect 884 30 890 32
<< pdif >>
rect 77 363 82 375
rect 75 361 82 363
rect 75 359 77 361
rect 79 359 82 361
rect 75 354 82 359
rect 75 352 77 354
rect 79 352 82 354
rect 75 350 82 352
rect 84 373 93 375
rect 84 371 88 373
rect 90 371 93 373
rect 116 373 130 375
rect 116 372 123 373
rect 84 363 93 371
rect 100 363 105 372
rect 84 350 95 363
rect 97 354 105 363
rect 97 352 100 354
rect 102 352 105 354
rect 97 350 105 352
rect 100 347 105 350
rect 107 347 112 372
rect 114 371 123 372
rect 125 371 130 373
rect 114 366 130 371
rect 114 364 123 366
rect 125 364 130 366
rect 114 347 130 364
rect 132 365 140 375
rect 132 363 135 365
rect 137 363 140 365
rect 132 358 140 363
rect 132 356 135 358
rect 137 356 140 358
rect 132 347 140 356
rect 142 373 150 375
rect 142 371 145 373
rect 147 371 150 373
rect 142 366 150 371
rect 142 364 145 366
rect 147 364 150 366
rect 142 347 150 364
rect 152 360 157 375
rect 177 363 182 375
rect 175 361 182 363
rect 152 358 159 360
rect 152 356 155 358
rect 157 356 159 358
rect 152 351 159 356
rect 152 349 155 351
rect 157 349 159 351
rect 175 359 177 361
rect 179 359 182 361
rect 175 354 182 359
rect 175 352 177 354
rect 179 352 182 354
rect 175 350 182 352
rect 184 373 193 375
rect 184 371 188 373
rect 190 371 193 373
rect 216 373 230 375
rect 216 372 223 373
rect 184 363 193 371
rect 200 363 205 372
rect 184 350 195 363
rect 197 354 205 363
rect 197 352 200 354
rect 202 352 205 354
rect 197 350 205 352
rect 152 347 159 349
rect 200 347 205 350
rect 207 347 212 372
rect 214 371 223 372
rect 225 371 230 373
rect 214 366 230 371
rect 214 364 223 366
rect 225 364 230 366
rect 214 347 230 364
rect 232 365 240 375
rect 232 363 235 365
rect 237 363 240 365
rect 232 358 240 363
rect 232 356 235 358
rect 237 356 240 358
rect 232 347 240 356
rect 242 373 250 375
rect 242 371 245 373
rect 247 371 250 373
rect 242 366 250 371
rect 242 364 245 366
rect 247 364 250 366
rect 242 347 250 364
rect 252 360 257 375
rect 275 373 284 375
rect 275 371 278 373
rect 280 371 284 373
rect 275 366 284 371
rect 264 364 271 366
rect 264 362 266 364
rect 268 362 271 364
rect 264 360 271 362
rect 252 358 259 360
rect 252 356 255 358
rect 257 356 259 358
rect 252 351 259 356
rect 266 354 271 360
rect 273 357 284 366
rect 286 357 291 375
rect 293 368 298 375
rect 293 366 300 368
rect 293 364 296 366
rect 298 364 300 366
rect 293 362 300 364
rect 306 363 311 375
rect 293 357 298 362
rect 304 361 311 363
rect 304 359 306 361
rect 308 359 311 361
rect 273 354 281 357
rect 252 349 255 351
rect 257 349 259 351
rect 252 347 259 349
rect 304 354 311 359
rect 304 352 306 354
rect 308 352 311 354
rect 304 350 311 352
rect 313 373 322 375
rect 313 371 317 373
rect 319 371 322 373
rect 345 373 359 375
rect 345 372 352 373
rect 313 363 322 371
rect 329 363 334 372
rect 313 350 324 363
rect 326 354 334 363
rect 326 352 329 354
rect 331 352 334 354
rect 326 350 334 352
rect 329 347 334 350
rect 336 347 341 372
rect 343 371 352 372
rect 354 371 359 373
rect 343 366 359 371
rect 343 364 352 366
rect 354 364 359 366
rect 343 347 359 364
rect 361 365 369 375
rect 361 363 364 365
rect 366 363 369 365
rect 361 358 369 363
rect 361 356 364 358
rect 366 356 369 358
rect 361 347 369 356
rect 371 373 379 375
rect 371 371 374 373
rect 376 371 379 373
rect 371 366 379 371
rect 371 364 374 366
rect 376 364 379 366
rect 371 347 379 364
rect 381 360 386 375
rect 401 363 406 375
rect 399 361 406 363
rect 381 358 388 360
rect 381 356 384 358
rect 386 356 388 358
rect 381 351 388 356
rect 381 349 384 351
rect 386 349 388 351
rect 399 359 401 361
rect 403 359 406 361
rect 399 354 406 359
rect 399 352 401 354
rect 403 352 406 354
rect 399 350 406 352
rect 408 373 417 375
rect 408 371 412 373
rect 414 371 417 373
rect 440 373 454 375
rect 440 372 447 373
rect 408 363 417 371
rect 424 363 429 372
rect 408 350 419 363
rect 421 354 429 363
rect 421 352 424 354
rect 426 352 429 354
rect 421 350 429 352
rect 381 347 388 349
rect 424 347 429 350
rect 431 347 436 372
rect 438 371 447 372
rect 449 371 454 373
rect 438 366 454 371
rect 438 364 447 366
rect 449 364 454 366
rect 438 347 454 364
rect 456 365 464 375
rect 456 363 459 365
rect 461 363 464 365
rect 456 358 464 363
rect 456 356 459 358
rect 461 356 464 358
rect 456 347 464 356
rect 466 373 474 375
rect 466 371 469 373
rect 471 371 474 373
rect 466 366 474 371
rect 466 364 469 366
rect 471 364 474 366
rect 466 347 474 364
rect 476 360 481 375
rect 499 373 508 375
rect 499 371 502 373
rect 504 371 508 373
rect 499 366 508 371
rect 488 364 495 366
rect 488 362 490 364
rect 492 362 495 364
rect 488 360 495 362
rect 476 358 483 360
rect 476 356 479 358
rect 481 356 483 358
rect 476 351 483 356
rect 490 354 495 360
rect 497 357 508 366
rect 510 357 515 375
rect 517 368 522 375
rect 517 366 524 368
rect 517 364 520 366
rect 522 364 524 366
rect 517 362 524 364
rect 530 363 535 375
rect 517 357 522 362
rect 528 361 535 363
rect 528 359 530 361
rect 532 359 535 361
rect 497 354 505 357
rect 476 349 479 351
rect 481 349 483 351
rect 476 347 483 349
rect 528 354 535 359
rect 528 352 530 354
rect 532 352 535 354
rect 528 350 535 352
rect 537 373 546 375
rect 537 371 541 373
rect 543 371 546 373
rect 569 373 583 375
rect 569 372 576 373
rect 537 363 546 371
rect 553 363 558 372
rect 537 350 548 363
rect 550 354 558 363
rect 550 352 553 354
rect 555 352 558 354
rect 550 350 558 352
rect 553 347 558 350
rect 560 347 565 372
rect 567 371 576 372
rect 578 371 583 373
rect 567 366 583 371
rect 567 364 576 366
rect 578 364 583 366
rect 567 347 583 364
rect 585 365 593 375
rect 585 363 588 365
rect 590 363 593 365
rect 585 358 593 363
rect 585 356 588 358
rect 590 356 593 358
rect 585 347 593 356
rect 595 373 603 375
rect 595 371 598 373
rect 600 371 603 373
rect 595 366 603 371
rect 595 364 598 366
rect 600 364 603 366
rect 595 347 603 364
rect 605 360 610 375
rect 626 363 631 375
rect 624 361 631 363
rect 605 358 612 360
rect 605 356 608 358
rect 610 356 612 358
rect 605 351 612 356
rect 605 349 608 351
rect 610 349 612 351
rect 624 359 626 361
rect 628 359 631 361
rect 624 354 631 359
rect 624 352 626 354
rect 628 352 631 354
rect 624 350 631 352
rect 633 373 642 375
rect 633 371 637 373
rect 639 371 642 373
rect 665 373 679 375
rect 665 372 672 373
rect 633 363 642 371
rect 649 363 654 372
rect 633 350 644 363
rect 646 354 654 363
rect 646 352 649 354
rect 651 352 654 354
rect 646 350 654 352
rect 605 347 612 349
rect 649 347 654 350
rect 656 347 661 372
rect 663 371 672 372
rect 674 371 679 373
rect 663 366 679 371
rect 663 364 672 366
rect 674 364 679 366
rect 663 347 679 364
rect 681 365 689 375
rect 681 363 684 365
rect 686 363 689 365
rect 681 358 689 363
rect 681 356 684 358
rect 686 356 689 358
rect 681 347 689 356
rect 691 373 699 375
rect 691 371 694 373
rect 696 371 699 373
rect 691 366 699 371
rect 691 364 694 366
rect 696 364 699 366
rect 691 347 699 364
rect 701 360 706 375
rect 701 358 708 360
rect 701 356 704 358
rect 706 356 708 358
rect 701 351 708 356
rect 725 353 730 359
rect 701 349 704 351
rect 706 349 708 351
rect 701 347 708 349
rect 723 351 730 353
rect 723 349 725 351
rect 727 349 730 351
rect 723 347 730 349
rect 732 357 738 359
rect 732 351 740 357
rect 732 349 735 351
rect 737 349 740 351
rect 732 347 740 349
rect 742 351 750 357
rect 742 349 745 351
rect 747 349 750 351
rect 742 347 750 349
rect 752 355 759 357
rect 752 353 755 355
rect 757 353 759 355
rect 774 353 779 359
rect 752 347 759 353
rect 772 351 779 353
rect 772 349 774 351
rect 776 349 779 351
rect 772 347 779 349
rect 781 357 787 359
rect 781 351 789 357
rect 781 349 784 351
rect 786 349 789 351
rect 781 347 789 349
rect 791 351 799 357
rect 791 349 794 351
rect 796 349 799 351
rect 791 347 799 349
rect 801 355 808 357
rect 801 353 804 355
rect 806 353 808 355
rect 824 353 829 359
rect 801 347 808 353
rect 822 351 829 353
rect 822 349 824 351
rect 826 349 829 351
rect 822 347 829 349
rect 831 357 837 359
rect 831 351 839 357
rect 831 349 834 351
rect 836 349 839 351
rect 831 347 839 349
rect 841 351 849 357
rect 841 349 844 351
rect 846 349 849 351
rect 841 347 849 349
rect 851 355 858 357
rect 851 353 854 355
rect 856 353 858 355
rect 851 347 858 353
rect 77 259 82 265
rect 75 257 82 259
rect 75 255 77 257
rect 79 255 82 257
rect 75 253 82 255
rect 84 263 90 265
rect 84 257 92 263
rect 84 255 87 257
rect 89 255 92 257
rect 84 253 92 255
rect 94 257 102 263
rect 94 255 97 257
rect 99 255 102 257
rect 94 253 102 255
rect 104 261 111 263
rect 104 259 107 261
rect 109 259 111 261
rect 127 259 132 265
rect 104 253 111 259
rect 125 257 132 259
rect 125 255 127 257
rect 129 255 132 257
rect 125 253 132 255
rect 134 263 140 265
rect 134 257 142 263
rect 134 255 137 257
rect 139 255 142 257
rect 134 253 142 255
rect 144 257 152 263
rect 144 255 147 257
rect 149 255 152 257
rect 144 253 152 255
rect 154 261 161 263
rect 154 259 157 261
rect 159 259 161 261
rect 198 260 203 266
rect 154 253 161 259
rect 196 258 203 260
rect 196 256 198 258
rect 200 256 203 258
rect 196 254 203 256
rect 205 264 211 266
rect 205 258 213 264
rect 205 256 208 258
rect 210 256 213 258
rect 205 254 213 256
rect 215 258 223 264
rect 215 256 218 258
rect 220 256 223 258
rect 215 254 223 256
rect 225 262 232 264
rect 225 260 228 262
rect 230 260 232 262
rect 239 260 244 266
rect 225 254 232 260
rect 237 258 244 260
rect 237 256 239 258
rect 241 256 244 258
rect 237 254 244 256
rect 246 264 252 266
rect 246 258 254 264
rect 246 256 249 258
rect 251 256 254 258
rect 246 254 254 256
rect 256 258 264 264
rect 256 256 259 258
rect 261 256 264 258
rect 256 254 264 256
rect 266 262 273 264
rect 266 260 269 262
rect 271 260 273 262
rect 266 254 273 260
rect 327 259 332 265
rect 325 257 332 259
rect 325 255 327 257
rect 329 255 332 257
rect 325 253 332 255
rect 334 263 340 265
rect 334 257 342 263
rect 334 255 337 257
rect 339 255 342 257
rect 334 253 342 255
rect 344 257 352 263
rect 344 255 347 257
rect 349 255 352 257
rect 344 253 352 255
rect 354 261 361 263
rect 354 259 357 261
rect 359 259 361 261
rect 377 259 382 265
rect 354 253 361 259
rect 375 257 382 259
rect 375 255 377 257
rect 379 255 382 257
rect 375 253 382 255
rect 384 263 390 265
rect 384 257 392 263
rect 384 255 387 257
rect 389 255 392 257
rect 384 253 392 255
rect 394 257 402 263
rect 394 255 397 257
rect 399 255 402 257
rect 394 253 402 255
rect 404 261 411 263
rect 404 259 407 261
rect 409 259 411 261
rect 421 259 426 265
rect 404 253 411 259
rect 419 257 426 259
rect 419 255 421 257
rect 423 255 426 257
rect 419 253 426 255
rect 428 263 434 265
rect 428 257 436 263
rect 428 255 431 257
rect 433 255 436 257
rect 428 253 436 255
rect 438 257 446 263
rect 438 255 441 257
rect 443 255 446 257
rect 438 253 446 255
rect 448 261 455 263
rect 448 259 451 261
rect 453 259 455 261
rect 477 259 482 265
rect 448 253 455 259
rect 475 257 482 259
rect 475 255 477 257
rect 479 255 482 257
rect 475 253 482 255
rect 484 263 490 265
rect 484 257 492 263
rect 484 255 487 257
rect 489 255 492 257
rect 484 253 492 255
rect 494 257 502 263
rect 494 255 497 257
rect 499 255 502 257
rect 494 253 502 255
rect 504 261 511 263
rect 504 259 507 261
rect 509 259 511 261
rect 527 259 532 265
rect 504 253 511 259
rect 525 257 532 259
rect 525 255 527 257
rect 529 255 532 257
rect 525 253 532 255
rect 534 263 540 265
rect 534 257 542 263
rect 534 255 537 257
rect 539 255 542 257
rect 534 253 542 255
rect 544 257 552 263
rect 544 255 547 257
rect 549 255 552 257
rect 544 253 552 255
rect 554 261 561 263
rect 554 259 557 261
rect 559 259 561 261
rect 577 259 582 265
rect 554 253 561 259
rect 575 257 582 259
rect 575 255 577 257
rect 579 255 582 257
rect 575 253 582 255
rect 584 263 590 265
rect 671 269 676 281
rect 584 257 592 263
rect 584 255 587 257
rect 589 255 592 257
rect 584 253 592 255
rect 594 257 602 263
rect 594 255 597 257
rect 599 255 602 257
rect 594 253 602 255
rect 604 261 611 263
rect 604 259 607 261
rect 609 259 611 261
rect 627 259 632 265
rect 604 253 611 259
rect 625 257 632 259
rect 625 255 627 257
rect 629 255 632 257
rect 625 253 632 255
rect 634 263 640 265
rect 669 267 676 269
rect 669 265 671 267
rect 673 265 676 267
rect 634 257 642 263
rect 634 255 637 257
rect 639 255 642 257
rect 634 253 642 255
rect 644 257 652 263
rect 644 255 647 257
rect 649 255 652 257
rect 644 253 652 255
rect 654 261 661 263
rect 654 259 657 261
rect 659 259 661 261
rect 654 253 661 259
rect 669 260 676 265
rect 669 258 671 260
rect 673 258 676 260
rect 669 256 676 258
rect 678 279 687 281
rect 678 277 682 279
rect 684 277 687 279
rect 710 279 724 281
rect 710 278 717 279
rect 678 269 687 277
rect 694 269 699 278
rect 678 256 689 269
rect 691 260 699 269
rect 691 258 694 260
rect 696 258 699 260
rect 691 256 699 258
rect 694 253 699 256
rect 701 253 706 278
rect 708 277 717 278
rect 719 277 724 279
rect 708 272 724 277
rect 708 270 717 272
rect 719 270 724 272
rect 708 253 724 270
rect 726 271 734 281
rect 726 269 729 271
rect 731 269 734 271
rect 726 264 734 269
rect 726 262 729 264
rect 731 262 734 264
rect 726 253 734 262
rect 736 279 744 281
rect 736 277 739 279
rect 741 277 744 279
rect 736 272 744 277
rect 736 270 739 272
rect 741 270 744 272
rect 736 253 744 270
rect 746 266 751 281
rect 771 269 776 281
rect 769 267 776 269
rect 746 264 753 266
rect 746 262 749 264
rect 751 262 753 264
rect 746 257 753 262
rect 746 255 749 257
rect 751 255 753 257
rect 769 265 771 267
rect 773 265 776 267
rect 769 260 776 265
rect 769 258 771 260
rect 773 258 776 260
rect 769 256 776 258
rect 778 279 787 281
rect 778 277 782 279
rect 784 277 787 279
rect 810 279 824 281
rect 810 278 817 279
rect 778 269 787 277
rect 794 269 799 278
rect 778 256 789 269
rect 791 260 799 269
rect 791 258 794 260
rect 796 258 799 260
rect 791 256 799 258
rect 746 253 753 255
rect 794 253 799 256
rect 801 253 806 278
rect 808 277 817 278
rect 819 277 824 279
rect 808 272 824 277
rect 808 270 817 272
rect 819 270 824 272
rect 808 253 824 270
rect 826 271 834 281
rect 826 269 829 271
rect 831 269 834 271
rect 826 264 834 269
rect 826 262 829 264
rect 831 262 834 264
rect 826 253 834 262
rect 836 279 844 281
rect 836 277 839 279
rect 841 277 844 279
rect 836 272 844 277
rect 836 270 839 272
rect 841 270 844 272
rect 836 253 844 270
rect 846 266 851 281
rect 846 264 853 266
rect 846 262 849 264
rect 851 262 853 264
rect 846 257 853 262
rect 846 255 849 257
rect 851 255 853 257
rect 846 253 853 255
rect 77 175 82 187
rect 75 173 82 175
rect 75 171 77 173
rect 79 171 82 173
rect 75 166 82 171
rect 75 164 77 166
rect 79 164 82 166
rect 75 162 82 164
rect 84 185 93 187
rect 84 183 88 185
rect 90 183 93 185
rect 116 185 130 187
rect 116 184 123 185
rect 84 175 93 183
rect 100 175 105 184
rect 84 162 95 175
rect 97 166 105 175
rect 97 164 100 166
rect 102 164 105 166
rect 97 162 105 164
rect 100 159 105 162
rect 107 159 112 184
rect 114 183 123 184
rect 125 183 130 185
rect 114 178 130 183
rect 114 176 123 178
rect 125 176 130 178
rect 114 159 130 176
rect 132 177 140 187
rect 132 175 135 177
rect 137 175 140 177
rect 132 170 140 175
rect 132 168 135 170
rect 137 168 140 170
rect 132 159 140 168
rect 142 185 150 187
rect 142 183 145 185
rect 147 183 150 185
rect 142 178 150 183
rect 142 176 145 178
rect 147 176 150 178
rect 142 159 150 176
rect 152 172 157 187
rect 175 185 184 187
rect 175 183 178 185
rect 180 183 184 185
rect 175 178 184 183
rect 164 176 171 178
rect 164 174 166 176
rect 168 174 171 176
rect 164 172 171 174
rect 152 170 159 172
rect 152 168 155 170
rect 157 168 159 170
rect 152 163 159 168
rect 166 166 171 172
rect 173 169 184 178
rect 186 169 191 187
rect 193 180 198 187
rect 193 178 200 180
rect 193 176 196 178
rect 198 176 200 178
rect 193 174 200 176
rect 206 175 211 187
rect 193 169 198 174
rect 204 173 211 175
rect 204 171 206 173
rect 208 171 211 173
rect 173 166 181 169
rect 152 161 155 163
rect 157 161 159 163
rect 152 159 159 161
rect 204 166 211 171
rect 204 164 206 166
rect 208 164 211 166
rect 204 162 211 164
rect 213 185 222 187
rect 213 183 217 185
rect 219 183 222 185
rect 245 185 259 187
rect 245 184 252 185
rect 213 175 222 183
rect 229 175 234 184
rect 213 162 224 175
rect 226 166 234 175
rect 226 164 229 166
rect 231 164 234 166
rect 226 162 234 164
rect 229 159 234 162
rect 236 159 241 184
rect 243 183 252 184
rect 254 183 259 185
rect 243 178 259 183
rect 243 176 252 178
rect 254 176 259 178
rect 243 159 259 176
rect 261 177 269 187
rect 261 175 264 177
rect 266 175 269 177
rect 261 170 269 175
rect 261 168 264 170
rect 266 168 269 170
rect 261 159 269 168
rect 271 185 279 187
rect 271 183 274 185
rect 276 183 279 185
rect 271 178 279 183
rect 271 176 274 178
rect 276 176 279 178
rect 271 159 279 176
rect 281 172 286 187
rect 301 175 306 187
rect 299 173 306 175
rect 281 170 288 172
rect 281 168 284 170
rect 286 168 288 170
rect 281 163 288 168
rect 281 161 284 163
rect 286 161 288 163
rect 299 171 301 173
rect 303 171 306 173
rect 299 166 306 171
rect 299 164 301 166
rect 303 164 306 166
rect 299 162 306 164
rect 308 185 317 187
rect 308 183 312 185
rect 314 183 317 185
rect 340 185 354 187
rect 340 184 347 185
rect 308 175 317 183
rect 324 175 329 184
rect 308 162 319 175
rect 321 166 329 175
rect 321 164 324 166
rect 326 164 329 166
rect 321 162 329 164
rect 281 159 288 161
rect 324 159 329 162
rect 331 159 336 184
rect 338 183 347 184
rect 349 183 354 185
rect 338 178 354 183
rect 338 176 347 178
rect 349 176 354 178
rect 338 159 354 176
rect 356 177 364 187
rect 356 175 359 177
rect 361 175 364 177
rect 356 170 364 175
rect 356 168 359 170
rect 361 168 364 170
rect 356 159 364 168
rect 366 185 374 187
rect 366 183 369 185
rect 371 183 374 185
rect 366 178 374 183
rect 366 176 369 178
rect 371 176 374 178
rect 366 159 374 176
rect 376 172 381 187
rect 399 185 408 187
rect 399 183 402 185
rect 404 183 408 185
rect 399 178 408 183
rect 388 176 395 178
rect 388 174 390 176
rect 392 174 395 176
rect 388 172 395 174
rect 376 170 383 172
rect 376 168 379 170
rect 381 168 383 170
rect 376 163 383 168
rect 390 166 395 172
rect 397 169 408 178
rect 410 169 415 187
rect 417 180 422 187
rect 417 178 424 180
rect 417 176 420 178
rect 422 176 424 178
rect 417 174 424 176
rect 430 175 435 187
rect 417 169 422 174
rect 428 173 435 175
rect 428 171 430 173
rect 432 171 435 173
rect 397 166 405 169
rect 376 161 379 163
rect 381 161 383 163
rect 376 159 383 161
rect 428 166 435 171
rect 428 164 430 166
rect 432 164 435 166
rect 428 162 435 164
rect 437 185 446 187
rect 437 183 441 185
rect 443 183 446 185
rect 469 185 483 187
rect 469 184 476 185
rect 437 175 446 183
rect 453 175 458 184
rect 437 162 448 175
rect 450 166 458 175
rect 450 164 453 166
rect 455 164 458 166
rect 450 162 458 164
rect 453 159 458 162
rect 460 159 465 184
rect 467 183 476 184
rect 478 183 483 185
rect 467 178 483 183
rect 467 176 476 178
rect 478 176 483 178
rect 467 159 483 176
rect 485 177 493 187
rect 485 175 488 177
rect 490 175 493 177
rect 485 170 493 175
rect 485 168 488 170
rect 490 168 493 170
rect 485 159 493 168
rect 495 185 503 187
rect 495 183 498 185
rect 500 183 503 185
rect 495 178 503 183
rect 495 176 498 178
rect 500 176 503 178
rect 495 159 503 176
rect 505 172 510 187
rect 525 175 530 187
rect 523 173 530 175
rect 505 170 512 172
rect 505 168 508 170
rect 510 168 512 170
rect 505 163 512 168
rect 505 161 508 163
rect 510 161 512 163
rect 523 171 525 173
rect 527 171 530 173
rect 523 166 530 171
rect 523 164 525 166
rect 527 164 530 166
rect 523 162 530 164
rect 532 185 541 187
rect 532 183 536 185
rect 538 183 541 185
rect 564 185 578 187
rect 564 184 571 185
rect 532 175 541 183
rect 548 175 553 184
rect 532 162 543 175
rect 545 166 553 175
rect 545 164 548 166
rect 550 164 553 166
rect 545 162 553 164
rect 505 159 512 161
rect 548 159 553 162
rect 555 159 560 184
rect 562 183 571 184
rect 573 183 578 185
rect 562 178 578 183
rect 562 176 571 178
rect 573 176 578 178
rect 562 159 578 176
rect 580 177 588 187
rect 580 175 583 177
rect 585 175 588 177
rect 580 170 588 175
rect 580 168 583 170
rect 585 168 588 170
rect 580 159 588 168
rect 590 185 598 187
rect 590 183 593 185
rect 595 183 598 185
rect 590 178 598 183
rect 590 176 593 178
rect 595 176 598 178
rect 590 159 598 176
rect 600 172 605 187
rect 623 185 632 187
rect 623 183 626 185
rect 628 183 632 185
rect 623 178 632 183
rect 612 176 619 178
rect 612 174 614 176
rect 616 174 619 176
rect 612 172 619 174
rect 600 170 607 172
rect 600 168 603 170
rect 605 168 607 170
rect 600 163 607 168
rect 614 166 619 172
rect 621 169 632 178
rect 634 169 639 187
rect 641 180 646 187
rect 641 178 648 180
rect 641 176 644 178
rect 646 176 648 178
rect 641 174 648 176
rect 654 175 659 187
rect 641 169 646 174
rect 652 173 659 175
rect 652 171 654 173
rect 656 171 659 173
rect 621 166 629 169
rect 600 161 603 163
rect 605 161 607 163
rect 600 159 607 161
rect 652 166 659 171
rect 652 164 654 166
rect 656 164 659 166
rect 652 162 659 164
rect 661 185 670 187
rect 661 183 665 185
rect 667 183 670 185
rect 693 185 707 187
rect 693 184 700 185
rect 661 175 670 183
rect 677 175 682 184
rect 661 162 672 175
rect 674 166 682 175
rect 674 164 677 166
rect 679 164 682 166
rect 674 162 682 164
rect 677 159 682 162
rect 684 159 689 184
rect 691 183 700 184
rect 702 183 707 185
rect 691 178 707 183
rect 691 176 700 178
rect 702 176 707 178
rect 691 159 707 176
rect 709 177 717 187
rect 709 175 712 177
rect 714 175 717 177
rect 709 170 717 175
rect 709 168 712 170
rect 714 168 717 170
rect 709 159 717 168
rect 719 185 727 187
rect 719 183 722 185
rect 724 183 727 185
rect 719 178 727 183
rect 719 176 722 178
rect 724 176 727 178
rect 719 159 727 176
rect 729 172 734 187
rect 729 170 736 172
rect 729 168 732 170
rect 734 168 736 170
rect 729 163 736 168
rect 749 165 754 171
rect 729 161 732 163
rect 734 161 736 163
rect 729 159 736 161
rect 747 163 754 165
rect 747 161 749 163
rect 751 161 754 163
rect 747 159 754 161
rect 756 169 762 171
rect 756 163 764 169
rect 756 161 759 163
rect 761 161 764 163
rect 756 159 764 161
rect 766 163 774 169
rect 766 161 769 163
rect 771 161 774 163
rect 766 159 774 161
rect 776 167 783 169
rect 776 165 779 167
rect 781 165 783 167
rect 776 159 783 165
rect 120 81 125 93
rect 76 71 81 77
rect 74 69 81 71
rect 74 67 76 69
rect 78 67 81 69
rect 74 65 81 67
rect 83 75 89 77
rect 118 79 125 81
rect 118 77 120 79
rect 122 77 125 79
rect 83 69 91 75
rect 83 67 86 69
rect 88 67 91 69
rect 83 65 91 67
rect 93 69 101 75
rect 93 67 96 69
rect 98 67 101 69
rect 93 65 101 67
rect 103 73 110 75
rect 103 71 106 73
rect 108 71 110 73
rect 103 65 110 71
rect 118 72 125 77
rect 118 70 120 72
rect 122 70 125 72
rect 118 68 125 70
rect 127 91 136 93
rect 127 89 131 91
rect 133 89 136 91
rect 159 91 173 93
rect 159 90 166 91
rect 127 81 136 89
rect 143 81 148 90
rect 127 68 138 81
rect 140 72 148 81
rect 140 70 143 72
rect 145 70 148 72
rect 140 68 148 70
rect 143 65 148 68
rect 150 65 155 90
rect 157 89 166 90
rect 168 89 173 91
rect 157 84 173 89
rect 157 82 166 84
rect 168 82 173 84
rect 157 65 173 82
rect 175 83 183 93
rect 175 81 178 83
rect 180 81 183 83
rect 175 76 183 81
rect 175 74 178 76
rect 180 74 183 76
rect 175 65 183 74
rect 185 91 193 93
rect 185 89 188 91
rect 190 89 193 91
rect 185 84 193 89
rect 185 82 188 84
rect 190 82 193 84
rect 185 65 193 82
rect 195 78 200 93
rect 218 91 227 93
rect 218 89 221 91
rect 223 89 227 91
rect 218 84 227 89
rect 207 82 214 84
rect 207 80 209 82
rect 211 80 214 82
rect 207 78 214 80
rect 195 76 202 78
rect 195 74 198 76
rect 200 74 202 76
rect 195 69 202 74
rect 209 72 214 78
rect 216 75 227 84
rect 229 75 234 93
rect 236 86 241 93
rect 236 84 243 86
rect 236 82 239 84
rect 241 82 243 84
rect 236 80 243 82
rect 249 81 254 93
rect 236 75 241 80
rect 247 79 254 81
rect 247 77 249 79
rect 251 77 254 79
rect 216 72 224 75
rect 195 67 198 69
rect 200 67 202 69
rect 195 65 202 67
rect 247 72 254 77
rect 247 70 249 72
rect 251 70 254 72
rect 247 68 254 70
rect 256 91 265 93
rect 256 89 260 91
rect 262 89 265 91
rect 288 91 302 93
rect 288 90 295 91
rect 256 81 265 89
rect 272 81 277 90
rect 256 68 267 81
rect 269 72 277 81
rect 269 70 272 72
rect 274 70 277 72
rect 269 68 277 70
rect 272 65 277 68
rect 279 65 284 90
rect 286 89 295 90
rect 297 89 302 91
rect 286 84 302 89
rect 286 82 295 84
rect 297 82 302 84
rect 286 65 302 82
rect 304 83 312 93
rect 304 81 307 83
rect 309 81 312 83
rect 304 76 312 81
rect 304 74 307 76
rect 309 74 312 76
rect 304 65 312 74
rect 314 91 322 93
rect 314 89 317 91
rect 319 89 322 91
rect 314 84 322 89
rect 314 82 317 84
rect 319 82 322 84
rect 314 65 322 82
rect 324 78 329 93
rect 324 76 331 78
rect 386 81 391 93
rect 324 74 327 76
rect 329 74 331 76
rect 324 69 331 74
rect 343 71 348 77
rect 324 67 327 69
rect 329 67 331 69
rect 324 65 331 67
rect 341 69 348 71
rect 341 67 343 69
rect 345 67 348 69
rect 341 65 348 67
rect 350 75 356 77
rect 384 79 391 81
rect 384 77 386 79
rect 388 77 391 79
rect 350 69 358 75
rect 350 67 353 69
rect 355 67 358 69
rect 350 65 358 67
rect 360 69 368 75
rect 360 67 363 69
rect 365 67 368 69
rect 360 65 368 67
rect 370 73 377 75
rect 370 71 373 73
rect 375 71 377 73
rect 370 65 377 71
rect 384 72 391 77
rect 384 70 386 72
rect 388 70 391 72
rect 384 68 391 70
rect 393 91 402 93
rect 393 89 397 91
rect 399 89 402 91
rect 425 91 439 93
rect 425 90 432 91
rect 393 81 402 89
rect 409 81 414 90
rect 393 68 404 81
rect 406 72 414 81
rect 406 70 409 72
rect 411 70 414 72
rect 406 68 414 70
rect 409 65 414 68
rect 416 65 421 90
rect 423 89 432 90
rect 434 89 439 91
rect 423 84 439 89
rect 423 82 432 84
rect 434 82 439 84
rect 423 65 439 82
rect 441 83 449 93
rect 441 81 444 83
rect 446 81 449 83
rect 441 76 449 81
rect 441 74 444 76
rect 446 74 449 76
rect 441 65 449 74
rect 451 91 459 93
rect 451 89 454 91
rect 456 89 459 91
rect 451 84 459 89
rect 451 82 454 84
rect 456 82 459 84
rect 451 65 459 82
rect 461 78 466 93
rect 484 91 493 93
rect 484 89 487 91
rect 489 89 493 91
rect 484 84 493 89
rect 473 82 480 84
rect 473 80 475 82
rect 477 80 480 82
rect 473 78 480 80
rect 461 76 468 78
rect 461 74 464 76
rect 466 74 468 76
rect 461 69 468 74
rect 475 72 480 78
rect 482 75 493 84
rect 495 75 500 93
rect 502 86 507 93
rect 502 84 509 86
rect 502 82 505 84
rect 507 82 509 84
rect 502 80 509 82
rect 515 81 520 93
rect 502 75 507 80
rect 513 79 520 81
rect 513 77 515 79
rect 517 77 520 79
rect 482 72 490 75
rect 461 67 464 69
rect 466 67 468 69
rect 461 65 468 67
rect 513 72 520 77
rect 513 70 515 72
rect 517 70 520 72
rect 513 68 520 70
rect 522 91 531 93
rect 522 89 526 91
rect 528 89 531 91
rect 554 91 568 93
rect 554 90 561 91
rect 522 81 531 89
rect 538 81 543 90
rect 522 68 533 81
rect 535 72 543 81
rect 535 70 538 72
rect 540 70 543 72
rect 535 68 543 70
rect 538 65 543 68
rect 545 65 550 90
rect 552 89 561 90
rect 563 89 568 91
rect 552 84 568 89
rect 552 82 561 84
rect 563 82 568 84
rect 552 65 568 82
rect 570 83 578 93
rect 570 81 573 83
rect 575 81 578 83
rect 570 76 578 81
rect 570 74 573 76
rect 575 74 578 76
rect 570 65 578 74
rect 580 91 588 93
rect 580 89 583 91
rect 585 89 588 91
rect 580 84 588 89
rect 580 82 583 84
rect 585 82 588 84
rect 580 65 588 82
rect 590 78 595 93
rect 590 76 597 78
rect 652 81 657 93
rect 590 74 593 76
rect 595 74 597 76
rect 590 69 597 74
rect 610 71 615 77
rect 590 67 593 69
rect 595 67 597 69
rect 590 65 597 67
rect 608 69 615 71
rect 608 67 610 69
rect 612 67 615 69
rect 608 65 615 67
rect 617 75 623 77
rect 650 79 657 81
rect 650 77 652 79
rect 654 77 657 79
rect 617 69 625 75
rect 617 67 620 69
rect 622 67 625 69
rect 617 65 625 67
rect 627 69 635 75
rect 627 67 630 69
rect 632 67 635 69
rect 627 65 635 67
rect 637 73 644 75
rect 637 71 640 73
rect 642 71 644 73
rect 637 65 644 71
rect 650 72 657 77
rect 650 70 652 72
rect 654 70 657 72
rect 650 68 657 70
rect 659 91 668 93
rect 659 89 663 91
rect 665 89 668 91
rect 691 91 705 93
rect 691 90 698 91
rect 659 81 668 89
rect 675 81 680 90
rect 659 68 670 81
rect 672 72 680 81
rect 672 70 675 72
rect 677 70 680 72
rect 672 68 680 70
rect 675 65 680 68
rect 682 65 687 90
rect 689 89 698 90
rect 700 89 705 91
rect 689 84 705 89
rect 689 82 698 84
rect 700 82 705 84
rect 689 65 705 82
rect 707 83 715 93
rect 707 81 710 83
rect 712 81 715 83
rect 707 76 715 81
rect 707 74 710 76
rect 712 74 715 76
rect 707 65 715 74
rect 717 91 725 93
rect 717 89 720 91
rect 722 89 725 91
rect 717 84 725 89
rect 717 82 720 84
rect 722 82 725 84
rect 717 65 725 82
rect 727 78 732 93
rect 750 91 759 93
rect 750 89 753 91
rect 755 89 759 91
rect 750 84 759 89
rect 739 82 746 84
rect 739 80 741 82
rect 743 80 746 82
rect 739 78 746 80
rect 727 76 734 78
rect 727 74 730 76
rect 732 74 734 76
rect 727 69 734 74
rect 741 72 746 78
rect 748 75 759 84
rect 761 75 766 93
rect 768 86 773 93
rect 768 84 775 86
rect 768 82 771 84
rect 773 82 775 84
rect 768 80 775 82
rect 781 81 786 93
rect 768 75 773 80
rect 779 79 786 81
rect 779 77 781 79
rect 783 77 786 79
rect 748 72 756 75
rect 727 67 730 69
rect 732 67 734 69
rect 727 65 734 67
rect 779 72 786 77
rect 779 70 781 72
rect 783 70 786 72
rect 779 68 786 70
rect 788 91 797 93
rect 788 89 792 91
rect 794 89 797 91
rect 820 91 834 93
rect 820 90 827 91
rect 788 81 797 89
rect 804 81 809 90
rect 788 68 799 81
rect 801 72 809 81
rect 801 70 804 72
rect 806 70 809 72
rect 801 68 809 70
rect 804 65 809 68
rect 811 65 816 90
rect 818 89 827 90
rect 829 89 834 91
rect 818 84 834 89
rect 818 82 827 84
rect 829 82 834 84
rect 818 65 834 82
rect 836 83 844 93
rect 836 81 839 83
rect 841 81 844 83
rect 836 76 844 81
rect 836 74 839 76
rect 841 74 844 76
rect 836 65 844 74
rect 846 91 854 93
rect 846 89 849 91
rect 851 89 854 91
rect 846 84 854 89
rect 846 82 849 84
rect 851 82 854 84
rect 846 65 854 82
rect 856 78 861 93
rect 856 76 863 78
rect 856 74 859 76
rect 861 74 863 76
rect 856 69 863 74
rect 875 71 880 77
rect 856 67 859 69
rect 861 67 863 69
rect 856 65 863 67
rect 873 69 880 71
rect 873 67 875 69
rect 877 67 880 69
rect 873 65 880 67
rect 882 75 888 77
rect 882 69 890 75
rect 882 67 885 69
rect 887 67 890 69
rect 882 65 890 67
rect 892 69 900 75
rect 892 67 895 69
rect 897 67 900 69
rect 892 65 900 67
rect 902 73 909 75
rect 902 71 905 73
rect 907 71 909 73
rect 902 65 909 71
<< alu1 >>
rect 32 381 195 382
rect 32 376 862 381
rect 32 374 267 376
rect 269 374 491 376
rect 493 374 726 376
rect 728 374 740 376
rect 742 374 754 376
rect 756 374 775 376
rect 777 374 789 376
rect 791 374 803 376
rect 805 374 825 376
rect 827 374 839 376
rect 841 374 853 376
rect 855 374 862 376
rect 32 373 862 374
rect 32 288 47 373
rect 75 363 88 367
rect 175 366 188 367
rect 175 364 176 366
rect 178 364 188 366
rect 175 363 188 364
rect 264 364 277 367
rect 75 361 80 363
rect 75 359 77 361
rect 79 359 80 361
rect 175 361 180 363
rect 75 354 80 359
rect 75 352 77 354
rect 79 352 80 354
rect 75 350 80 352
rect 75 343 79 350
rect 75 341 76 343
rect 78 341 79 343
rect 106 347 144 351
rect 75 328 79 341
rect 106 344 111 347
rect 103 342 111 344
rect 103 340 104 342
rect 106 340 111 342
rect 103 338 111 340
rect 121 342 136 343
rect 121 340 123 342
rect 125 340 130 342
rect 132 340 136 342
rect 121 339 136 340
rect 75 326 80 328
rect 123 333 127 339
rect 154 358 160 360
rect 154 356 155 358
rect 157 356 160 358
rect 154 351 160 356
rect 154 349 155 351
rect 157 349 160 351
rect 154 347 160 349
rect 123 331 124 333
rect 126 331 127 333
rect 123 330 127 331
rect 156 328 160 347
rect 175 359 177 361
rect 179 359 180 361
rect 264 362 266 364
rect 268 363 277 364
rect 304 363 317 367
rect 399 366 412 367
rect 399 364 407 366
rect 409 364 412 366
rect 399 363 412 364
rect 488 364 501 367
rect 175 354 180 359
rect 175 352 177 354
rect 179 352 180 354
rect 175 350 180 352
rect 175 328 179 350
rect 206 350 244 351
rect 206 348 234 350
rect 236 348 244 350
rect 206 347 244 348
rect 206 344 211 347
rect 203 342 211 344
rect 203 340 204 342
rect 206 340 211 342
rect 203 338 211 340
rect 221 342 236 343
rect 221 340 223 342
rect 225 340 230 342
rect 232 340 236 342
rect 221 339 236 340
rect 156 327 166 328
rect 75 324 77 326
rect 79 324 80 326
rect 75 322 80 324
rect 138 326 166 327
rect 138 324 155 326
rect 157 325 166 326
rect 157 324 162 325
rect 138 323 162 324
rect 164 323 166 325
rect 156 322 166 323
rect 175 326 180 328
rect 223 333 227 339
rect 254 358 260 360
rect 254 356 255 358
rect 257 356 260 358
rect 254 351 260 356
rect 254 349 255 351
rect 257 349 260 351
rect 254 347 260 349
rect 223 331 224 333
rect 226 331 227 333
rect 223 330 227 331
rect 256 327 260 347
rect 175 324 177 326
rect 179 324 180 326
rect 175 322 180 324
rect 238 326 260 327
rect 238 324 255 326
rect 257 324 260 326
rect 238 323 260 324
rect 264 342 268 362
rect 304 361 309 363
rect 264 340 265 342
rect 267 340 268 342
rect 264 330 268 340
rect 288 351 292 360
rect 304 359 306 361
rect 308 359 309 361
rect 399 361 404 363
rect 304 354 309 359
rect 304 352 306 354
rect 308 352 309 354
rect 279 350 292 351
rect 279 348 280 350
rect 282 348 283 350
rect 285 348 292 350
rect 279 347 292 348
rect 296 351 300 352
rect 296 349 297 351
rect 299 349 300 351
rect 296 343 300 349
rect 287 342 300 343
rect 287 340 293 342
rect 295 340 300 342
rect 287 339 300 340
rect 296 338 300 339
rect 304 350 309 352
rect 304 342 308 350
rect 304 340 305 342
rect 307 340 308 342
rect 335 347 373 351
rect 264 328 269 330
rect 264 326 266 328
rect 268 326 269 328
rect 264 322 269 326
rect 304 328 308 340
rect 335 344 340 347
rect 332 342 340 344
rect 332 340 333 342
rect 335 340 340 342
rect 332 338 340 340
rect 350 342 365 343
rect 350 340 352 342
rect 354 340 359 342
rect 361 340 365 342
rect 350 339 365 340
rect 304 326 309 328
rect 352 334 356 339
rect 383 358 389 360
rect 383 356 384 358
rect 386 356 389 358
rect 383 351 389 356
rect 383 349 384 351
rect 386 349 389 351
rect 383 347 389 349
rect 352 332 353 334
rect 355 332 356 334
rect 352 330 356 332
rect 385 327 389 347
rect 304 324 306 326
rect 308 324 309 326
rect 304 322 309 324
rect 367 326 389 327
rect 367 324 384 326
rect 386 324 389 326
rect 367 323 389 324
rect 399 359 401 361
rect 403 359 404 361
rect 488 362 490 364
rect 492 363 501 364
rect 528 363 541 367
rect 624 363 637 367
rect 399 354 404 359
rect 399 352 401 354
rect 403 352 404 354
rect 399 350 404 352
rect 399 328 403 350
rect 430 350 468 351
rect 430 348 458 350
rect 460 348 468 350
rect 430 347 468 348
rect 430 344 435 347
rect 427 342 435 344
rect 427 340 428 342
rect 430 340 435 342
rect 427 338 435 340
rect 445 342 460 343
rect 445 340 447 342
rect 449 340 454 342
rect 456 340 460 342
rect 445 339 460 340
rect 399 326 404 328
rect 447 333 451 339
rect 478 358 484 360
rect 478 356 479 358
rect 481 356 484 358
rect 478 351 484 356
rect 478 349 479 351
rect 481 349 484 351
rect 478 347 484 349
rect 447 331 448 333
rect 450 331 451 333
rect 447 330 451 331
rect 480 327 484 347
rect 399 324 401 326
rect 403 324 404 326
rect 399 322 404 324
rect 462 326 484 327
rect 462 324 479 326
rect 481 324 484 326
rect 462 323 484 324
rect 488 342 492 362
rect 528 361 533 363
rect 488 340 489 342
rect 491 340 492 342
rect 488 330 492 340
rect 512 351 516 360
rect 528 359 530 361
rect 532 359 533 361
rect 624 361 629 363
rect 528 354 533 359
rect 528 352 530 354
rect 532 352 533 354
rect 503 350 516 351
rect 503 348 504 350
rect 506 348 507 350
rect 509 348 516 350
rect 503 347 516 348
rect 520 351 524 352
rect 520 349 521 351
rect 523 349 524 351
rect 520 343 524 349
rect 511 342 524 343
rect 511 340 517 342
rect 519 340 524 342
rect 511 339 524 340
rect 520 338 524 339
rect 528 350 533 352
rect 528 342 532 350
rect 528 340 529 342
rect 531 340 532 342
rect 559 347 597 351
rect 488 328 493 330
rect 488 326 490 328
rect 492 326 493 328
rect 488 322 493 326
rect 528 328 532 340
rect 559 344 564 347
rect 556 342 564 344
rect 556 340 557 342
rect 559 340 561 342
rect 563 340 564 342
rect 556 338 564 340
rect 574 342 589 343
rect 574 340 576 342
rect 578 340 583 342
rect 585 340 589 342
rect 574 339 589 340
rect 528 326 533 328
rect 576 333 580 339
rect 607 358 613 360
rect 607 356 608 358
rect 610 356 613 358
rect 607 351 613 356
rect 607 349 608 351
rect 610 349 613 351
rect 607 347 613 349
rect 576 331 577 333
rect 579 331 580 333
rect 576 330 580 331
rect 609 327 613 347
rect 528 324 530 326
rect 532 324 533 326
rect 528 322 533 324
rect 591 326 613 327
rect 591 324 608 326
rect 610 324 613 326
rect 591 323 613 324
rect 624 359 626 361
rect 628 359 629 361
rect 624 354 629 359
rect 624 352 626 354
rect 628 352 629 354
rect 624 350 629 352
rect 624 328 628 350
rect 655 347 693 351
rect 655 344 660 347
rect 652 342 660 344
rect 652 340 653 342
rect 655 341 660 342
rect 655 340 656 341
rect 652 339 656 340
rect 658 339 660 341
rect 670 342 685 343
rect 670 340 672 342
rect 674 340 679 342
rect 681 340 685 342
rect 670 339 685 340
rect 652 338 660 339
rect 672 335 676 339
rect 703 358 709 360
rect 703 356 704 358
rect 706 356 709 358
rect 703 354 709 356
rect 703 352 705 354
rect 707 352 709 354
rect 703 351 709 352
rect 703 349 704 351
rect 706 349 709 351
rect 703 347 709 349
rect 624 326 629 328
rect 672 333 673 335
rect 675 333 676 335
rect 672 330 676 333
rect 705 327 709 347
rect 624 324 626 326
rect 628 324 629 326
rect 624 322 629 324
rect 687 326 709 327
rect 687 324 704 326
rect 706 324 709 326
rect 687 323 709 324
rect 723 351 727 360
rect 723 349 725 351
rect 723 336 727 349
rect 738 366 751 368
rect 738 364 742 366
rect 744 364 751 366
rect 738 362 751 364
rect 738 355 744 362
rect 772 351 776 360
rect 772 349 774 351
rect 723 334 724 336
rect 726 334 727 336
rect 723 328 727 334
rect 723 326 725 328
rect 727 326 735 328
rect 723 322 735 326
rect 755 335 759 344
rect 746 334 759 335
rect 746 332 751 334
rect 753 332 759 334
rect 746 330 759 332
rect 772 338 776 349
rect 787 366 800 368
rect 787 364 791 366
rect 793 364 800 366
rect 787 362 800 364
rect 787 355 793 362
rect 822 351 826 360
rect 822 349 824 351
rect 772 336 773 338
rect 775 336 776 338
rect 772 328 776 336
rect 772 326 774 328
rect 776 326 784 328
rect 772 322 784 326
rect 804 335 808 344
rect 795 334 808 335
rect 795 332 800 334
rect 802 332 808 334
rect 795 330 808 332
rect 822 337 826 349
rect 837 366 850 368
rect 837 364 841 366
rect 843 364 850 366
rect 837 362 850 364
rect 837 355 843 362
rect 822 335 823 337
rect 825 335 826 337
rect 822 328 826 335
rect 822 326 824 328
rect 826 326 834 328
rect 822 322 834 326
rect 854 335 858 344
rect 845 334 858 335
rect 845 332 850 334
rect 852 332 858 334
rect 845 330 858 332
rect 892 317 903 318
rect 71 313 154 317
rect 174 316 911 317
rect 174 314 267 316
rect 269 314 295 316
rect 297 314 491 316
rect 493 314 519 316
rect 521 314 726 316
rect 728 314 736 316
rect 738 314 775 316
rect 777 314 785 316
rect 787 314 825 316
rect 827 314 835 316
rect 837 314 911 316
rect 174 313 911 314
rect 71 310 911 313
rect 71 309 862 310
rect 154 307 187 309
rect 28 287 75 288
rect 112 287 125 288
rect 164 287 327 288
rect 361 287 374 288
rect 415 287 578 289
rect 28 283 867 287
rect 28 282 199 283
rect 28 280 78 282
rect 80 280 92 282
rect 94 280 106 282
rect 108 280 128 282
rect 130 280 142 282
rect 144 280 156 282
rect 158 281 199 282
rect 201 281 213 283
rect 215 281 227 283
rect 229 281 240 283
rect 242 281 254 283
rect 256 281 268 283
rect 270 282 867 283
rect 270 281 328 282
rect 158 280 328 281
rect 330 280 342 282
rect 344 280 356 282
rect 358 280 378 282
rect 380 280 392 282
rect 394 280 406 282
rect 408 280 422 282
rect 424 280 436 282
rect 438 280 450 282
rect 452 280 478 282
rect 480 280 492 282
rect 494 280 506 282
rect 508 280 528 282
rect 530 280 542 282
rect 544 280 556 282
rect 558 280 578 282
rect 580 280 592 282
rect 594 280 606 282
rect 608 280 628 282
rect 630 280 642 282
rect 644 280 656 282
rect 658 280 867 282
rect 28 279 115 280
rect 121 279 192 280
rect 28 193 47 279
rect 75 257 79 266
rect 75 255 77 257
rect 75 245 79 255
rect 90 272 103 274
rect 90 270 94 272
rect 96 270 103 272
rect 90 268 103 270
rect 90 261 96 268
rect 125 257 129 266
rect 125 255 127 257
rect 75 243 76 245
rect 78 243 79 245
rect 75 234 79 243
rect 75 232 77 234
rect 79 232 87 234
rect 75 228 87 232
rect 107 241 111 250
rect 98 240 111 241
rect 98 238 103 240
rect 105 238 111 240
rect 98 236 111 238
rect 125 247 129 255
rect 140 272 153 274
rect 140 270 144 272
rect 146 270 153 272
rect 140 268 153 270
rect 140 261 146 268
rect 196 258 200 267
rect 196 256 198 258
rect 125 245 126 247
rect 128 245 129 247
rect 125 234 129 245
rect 125 232 127 234
rect 129 232 137 234
rect 125 228 137 232
rect 157 241 161 250
rect 148 240 161 241
rect 148 238 153 240
rect 155 238 161 240
rect 148 236 161 238
rect 196 235 200 256
rect 211 273 224 275
rect 211 271 215 273
rect 217 271 224 273
rect 211 269 224 271
rect 211 262 217 269
rect 236 279 245 280
rect 237 258 241 267
rect 237 256 239 258
rect 196 233 198 235
rect 200 233 208 235
rect 196 229 208 233
rect 228 242 232 251
rect 219 241 232 242
rect 219 239 224 241
rect 226 239 232 241
rect 219 237 232 239
rect 237 235 241 256
rect 265 279 268 280
rect 252 273 265 275
rect 252 271 256 273
rect 258 271 265 273
rect 252 269 265 271
rect 252 262 258 269
rect 288 279 365 280
rect 371 279 459 280
rect 471 279 565 280
rect 571 279 867 280
rect 325 257 329 266
rect 325 255 327 257
rect 237 233 239 235
rect 241 233 249 235
rect 237 229 249 233
rect 269 242 273 251
rect 260 241 273 242
rect 260 239 265 241
rect 267 239 273 241
rect 260 237 273 239
rect 325 244 329 255
rect 340 272 353 274
rect 340 270 344 272
rect 346 270 353 272
rect 340 268 353 270
rect 340 261 346 268
rect 375 257 379 266
rect 375 255 377 257
rect 325 242 326 244
rect 328 242 329 244
rect 325 234 329 242
rect 325 232 327 234
rect 329 232 337 234
rect 325 228 337 232
rect 357 241 361 250
rect 348 240 361 241
rect 348 238 353 240
rect 355 238 361 240
rect 348 236 361 238
rect 375 247 379 255
rect 390 272 403 274
rect 390 270 394 272
rect 396 270 403 272
rect 390 268 403 270
rect 390 261 396 268
rect 419 257 423 266
rect 419 255 421 257
rect 375 245 376 247
rect 378 245 379 247
rect 375 234 379 245
rect 375 232 377 234
rect 379 232 387 234
rect 375 228 387 232
rect 407 241 411 250
rect 398 240 411 241
rect 398 238 403 240
rect 405 238 411 240
rect 398 236 411 238
rect 419 234 423 255
rect 434 272 447 274
rect 434 270 438 272
rect 440 270 447 272
rect 434 268 447 270
rect 434 261 440 268
rect 475 257 479 266
rect 475 255 477 257
rect 419 232 421 234
rect 423 232 431 234
rect 419 228 431 232
rect 451 241 455 250
rect 442 240 455 241
rect 442 238 447 240
rect 449 238 455 240
rect 442 236 455 238
rect 475 241 479 255
rect 490 272 498 274
rect 490 270 494 272
rect 496 270 498 272
rect 490 268 498 270
rect 490 261 496 268
rect 525 257 529 266
rect 525 255 527 257
rect 475 239 476 241
rect 478 239 479 241
rect 475 234 479 239
rect 475 232 477 234
rect 479 232 487 234
rect 475 228 487 232
rect 507 241 511 250
rect 498 240 511 241
rect 498 238 503 240
rect 505 238 511 240
rect 498 236 511 238
rect 525 243 529 255
rect 540 272 553 274
rect 540 270 544 272
rect 546 270 553 272
rect 540 268 553 270
rect 540 261 546 268
rect 575 257 579 266
rect 575 255 577 257
rect 525 241 526 243
rect 528 241 529 243
rect 525 234 529 241
rect 525 232 527 234
rect 529 232 537 234
rect 525 228 537 232
rect 557 241 561 250
rect 548 240 561 241
rect 548 238 553 240
rect 555 238 561 240
rect 548 236 561 238
rect 575 244 579 255
rect 590 272 598 274
rect 590 270 594 272
rect 596 270 598 272
rect 590 268 598 270
rect 590 261 596 268
rect 625 257 629 266
rect 625 255 627 257
rect 575 242 576 244
rect 578 242 579 244
rect 575 234 579 242
rect 575 232 577 234
rect 579 232 587 234
rect 575 228 587 232
rect 607 241 611 250
rect 598 240 611 241
rect 598 238 603 240
rect 605 238 611 240
rect 598 236 611 238
rect 625 246 629 255
rect 640 272 653 274
rect 640 270 644 272
rect 646 270 650 272
rect 652 270 653 272
rect 640 268 653 270
rect 640 261 646 268
rect 669 269 682 273
rect 769 269 782 273
rect 669 267 674 269
rect 669 265 671 267
rect 673 265 674 267
rect 769 267 774 269
rect 669 260 674 265
rect 669 258 671 260
rect 673 258 674 260
rect 669 256 674 258
rect 625 244 626 246
rect 628 244 629 246
rect 625 234 629 244
rect 625 232 627 234
rect 629 232 637 234
rect 625 228 637 232
rect 657 241 661 250
rect 648 240 661 241
rect 648 238 653 240
rect 655 238 661 240
rect 648 236 661 238
rect 669 234 673 256
rect 700 253 738 257
rect 700 250 705 253
rect 697 248 705 250
rect 697 246 698 248
rect 700 246 701 248
rect 703 246 705 248
rect 697 244 705 246
rect 715 248 730 249
rect 715 246 717 248
rect 719 246 724 248
rect 726 246 730 248
rect 715 245 730 246
rect 669 232 674 234
rect 717 236 721 245
rect 748 264 754 266
rect 748 262 749 264
rect 751 262 754 264
rect 748 257 754 262
rect 748 255 749 257
rect 751 255 754 257
rect 748 253 754 255
rect 750 235 754 253
rect 748 233 754 235
rect 669 230 671 232
rect 673 230 674 232
rect 669 228 674 230
rect 732 232 754 233
rect 732 230 749 232
rect 751 230 754 232
rect 732 229 754 230
rect 769 265 771 267
rect 773 265 774 267
rect 769 260 774 265
rect 769 258 771 260
rect 773 258 774 260
rect 769 256 774 258
rect 769 234 773 256
rect 800 253 838 257
rect 800 250 805 253
rect 797 248 805 250
rect 797 246 798 248
rect 800 246 801 248
rect 803 246 805 248
rect 797 244 805 246
rect 815 248 830 249
rect 815 246 817 248
rect 819 246 824 248
rect 826 246 830 248
rect 815 245 830 246
rect 769 232 774 234
rect 817 239 821 245
rect 848 264 854 266
rect 848 262 849 264
rect 851 262 854 264
rect 848 257 854 262
rect 848 255 849 257
rect 851 255 854 257
rect 848 253 854 255
rect 817 237 818 239
rect 820 237 821 239
rect 817 236 821 237
rect 850 233 854 253
rect 769 230 771 232
rect 773 230 774 232
rect 769 228 774 230
rect 832 232 854 233
rect 832 230 849 232
rect 851 230 854 232
rect 832 229 854 230
rect 192 223 277 224
rect 892 223 903 310
rect 71 222 165 223
rect 192 222 199 223
rect 71 220 78 222
rect 80 220 88 222
rect 90 220 128 222
rect 130 220 138 222
rect 140 221 199 222
rect 201 221 209 223
rect 211 221 240 223
rect 242 221 250 223
rect 252 222 365 223
rect 371 222 515 223
rect 252 221 328 222
rect 140 220 328 221
rect 330 220 338 222
rect 340 220 378 222
rect 380 220 388 222
rect 390 220 422 222
rect 424 220 432 222
rect 434 220 478 222
rect 480 220 488 222
rect 490 221 515 222
rect 521 222 615 223
rect 521 221 528 222
rect 490 220 528 221
rect 530 220 538 222
rect 540 220 578 222
rect 580 220 588 222
rect 590 221 615 222
rect 621 222 905 223
rect 621 221 628 222
rect 590 220 628 221
rect 630 220 638 222
rect 640 220 905 222
rect 71 216 905 220
rect 71 215 218 216
rect 321 215 459 216
rect 471 215 867 216
rect 362 214 375 215
rect 511 213 524 215
rect 612 213 625 215
rect 28 188 786 193
rect 28 186 167 188
rect 169 186 391 188
rect 393 186 615 188
rect 617 186 750 188
rect 752 186 764 188
rect 766 186 778 188
rect 780 186 786 188
rect 28 185 786 186
rect 28 184 88 185
rect 90 184 114 185
rect 29 99 45 184
rect 75 175 88 179
rect 164 176 177 179
rect 75 173 80 175
rect 75 171 77 173
rect 79 171 80 173
rect 164 174 166 176
rect 168 175 177 176
rect 204 175 217 179
rect 299 175 312 179
rect 388 176 401 179
rect 75 166 80 171
rect 75 164 77 166
rect 79 164 80 166
rect 75 162 80 164
rect 75 157 79 162
rect 75 155 76 157
rect 78 155 79 157
rect 75 140 79 155
rect 106 159 144 163
rect 106 156 111 159
rect 103 154 111 156
rect 103 152 104 154
rect 106 152 111 154
rect 103 150 111 152
rect 121 154 136 155
rect 121 152 123 154
rect 125 152 130 154
rect 132 152 136 154
rect 121 151 136 152
rect 75 138 80 140
rect 123 145 127 151
rect 154 170 160 172
rect 154 168 155 170
rect 157 168 160 170
rect 154 163 160 168
rect 154 161 155 163
rect 157 161 160 163
rect 154 159 160 161
rect 123 143 124 145
rect 126 143 127 145
rect 123 142 127 143
rect 156 139 160 159
rect 75 136 77 138
rect 79 136 80 138
rect 75 134 80 136
rect 138 138 160 139
rect 138 136 155 138
rect 157 136 160 138
rect 138 135 160 136
rect 164 171 168 174
rect 204 173 209 175
rect 164 169 165 171
rect 167 169 168 171
rect 164 142 168 169
rect 188 163 192 172
rect 204 171 206 173
rect 208 171 209 173
rect 299 173 304 175
rect 204 166 209 171
rect 204 164 206 166
rect 208 164 209 166
rect 179 162 192 163
rect 179 160 180 162
rect 182 160 183 162
rect 185 160 192 162
rect 179 159 192 160
rect 196 163 200 164
rect 196 161 197 163
rect 199 161 200 163
rect 196 155 200 161
rect 187 154 200 155
rect 187 152 193 154
rect 195 152 200 154
rect 187 151 200 152
rect 196 150 200 151
rect 204 162 209 164
rect 204 154 208 162
rect 204 152 205 154
rect 207 152 208 154
rect 235 159 273 163
rect 164 140 169 142
rect 164 138 166 140
rect 168 138 169 140
rect 164 134 169 138
rect 204 140 208 152
rect 235 156 240 159
rect 232 154 240 156
rect 232 152 233 154
rect 235 152 240 154
rect 232 150 240 152
rect 250 154 265 155
rect 250 152 252 154
rect 254 152 259 154
rect 261 152 265 154
rect 250 151 265 152
rect 252 148 256 151
rect 283 170 289 172
rect 283 168 284 170
rect 286 168 289 170
rect 283 163 289 168
rect 283 161 284 163
rect 286 161 289 163
rect 283 159 289 161
rect 204 138 209 140
rect 252 146 253 148
rect 255 146 256 148
rect 252 142 256 146
rect 285 139 289 159
rect 299 171 301 173
rect 303 171 304 173
rect 388 174 390 176
rect 392 175 401 176
rect 428 175 441 179
rect 523 175 536 179
rect 612 176 625 179
rect 299 166 304 171
rect 299 164 301 166
rect 303 164 304 166
rect 299 162 304 164
rect 299 146 303 162
rect 330 159 368 163
rect 330 156 335 159
rect 327 154 335 156
rect 327 152 328 154
rect 330 152 335 154
rect 327 150 335 152
rect 345 154 360 155
rect 345 152 347 154
rect 349 152 354 154
rect 356 152 360 154
rect 345 151 360 152
rect 204 136 206 138
rect 208 136 209 138
rect 204 134 209 136
rect 267 138 289 139
rect 267 136 284 138
rect 286 136 289 138
rect 267 135 289 136
rect 298 143 303 146
rect 298 141 300 143
rect 302 141 303 143
rect 298 140 303 141
rect 298 134 304 140
rect 347 145 351 151
rect 378 170 384 172
rect 378 168 379 170
rect 381 168 384 170
rect 378 163 384 168
rect 378 161 379 163
rect 381 161 384 163
rect 378 159 384 161
rect 347 143 348 145
rect 350 143 351 145
rect 347 142 351 143
rect 380 139 384 159
rect 362 138 384 139
rect 362 136 379 138
rect 381 136 384 138
rect 362 135 384 136
rect 388 142 392 174
rect 428 173 433 175
rect 412 163 416 172
rect 428 171 430 173
rect 432 171 433 173
rect 523 173 528 175
rect 428 166 433 171
rect 428 164 430 166
rect 432 164 433 166
rect 403 162 416 163
rect 403 160 404 162
rect 406 160 407 162
rect 409 160 416 162
rect 403 159 416 160
rect 420 163 424 164
rect 420 161 421 163
rect 423 161 424 163
rect 420 155 424 161
rect 411 154 424 155
rect 411 152 417 154
rect 419 152 424 154
rect 411 151 424 152
rect 420 150 424 151
rect 428 162 433 164
rect 428 154 432 162
rect 428 152 429 154
rect 431 152 432 154
rect 459 159 497 163
rect 388 140 393 142
rect 388 138 390 140
rect 392 138 393 140
rect 388 134 393 138
rect 428 140 432 152
rect 459 156 464 159
rect 456 154 464 156
rect 456 152 457 154
rect 459 152 464 154
rect 456 150 464 152
rect 474 154 489 155
rect 474 152 476 154
rect 478 152 483 154
rect 485 152 489 154
rect 474 151 489 152
rect 476 148 480 151
rect 507 170 513 172
rect 507 168 508 170
rect 510 168 513 170
rect 507 163 513 168
rect 507 161 508 163
rect 510 161 513 163
rect 507 159 513 161
rect 428 138 433 140
rect 476 146 477 148
rect 479 146 480 148
rect 476 142 480 146
rect 509 139 513 159
rect 428 136 430 138
rect 432 136 433 138
rect 428 134 433 136
rect 491 138 513 139
rect 491 136 508 138
rect 510 136 513 138
rect 491 135 513 136
rect 523 171 525 173
rect 527 171 528 173
rect 612 174 614 176
rect 616 175 625 176
rect 652 175 665 179
rect 523 166 528 171
rect 523 164 525 166
rect 527 164 528 166
rect 523 162 528 164
rect 523 140 527 162
rect 554 159 592 163
rect 554 156 559 159
rect 551 154 559 156
rect 551 152 552 154
rect 554 152 559 154
rect 551 150 559 152
rect 569 154 584 155
rect 569 152 571 154
rect 573 152 578 154
rect 580 152 584 154
rect 569 151 584 152
rect 523 138 528 140
rect 571 145 575 151
rect 602 170 608 172
rect 602 168 603 170
rect 605 168 608 170
rect 602 163 608 168
rect 602 161 603 163
rect 605 161 608 163
rect 602 159 608 161
rect 571 143 572 145
rect 574 143 575 145
rect 571 142 575 143
rect 604 139 608 159
rect 523 136 525 138
rect 527 136 528 138
rect 523 134 528 136
rect 586 138 608 139
rect 586 136 603 138
rect 605 136 608 138
rect 586 135 608 136
rect 612 142 616 174
rect 652 173 657 175
rect 636 163 640 172
rect 652 171 654 173
rect 656 171 657 173
rect 652 166 657 171
rect 652 164 654 166
rect 656 164 657 166
rect 627 162 640 163
rect 627 160 628 162
rect 630 160 631 162
rect 633 160 640 162
rect 627 159 640 160
rect 644 163 648 164
rect 644 161 645 163
rect 647 161 648 163
rect 644 155 648 161
rect 635 154 648 155
rect 635 152 641 154
rect 643 152 648 154
rect 635 151 648 152
rect 644 150 648 151
rect 652 162 657 164
rect 652 154 656 162
rect 652 152 653 154
rect 655 152 656 154
rect 683 159 721 163
rect 612 140 617 142
rect 612 138 614 140
rect 616 138 617 140
rect 612 134 617 138
rect 652 140 656 152
rect 683 156 688 159
rect 680 154 688 156
rect 680 152 681 154
rect 683 152 688 154
rect 680 150 688 152
rect 698 154 713 155
rect 698 152 700 154
rect 702 152 707 154
rect 709 152 713 154
rect 698 151 713 152
rect 652 138 657 140
rect 700 146 704 151
rect 731 170 737 172
rect 731 168 732 170
rect 734 168 737 170
rect 731 163 737 168
rect 731 161 732 163
rect 734 161 737 163
rect 731 159 737 161
rect 700 144 701 146
rect 703 144 704 146
rect 700 142 704 144
rect 733 139 737 159
rect 652 136 654 138
rect 656 136 657 138
rect 652 134 657 136
rect 715 138 737 139
rect 715 136 732 138
rect 734 136 737 138
rect 715 135 737 136
rect 747 163 751 172
rect 747 161 749 163
rect 747 146 751 161
rect 762 178 775 180
rect 762 176 766 178
rect 768 176 775 178
rect 762 174 775 176
rect 762 167 768 174
rect 747 144 748 146
rect 750 144 751 146
rect 747 140 751 144
rect 747 138 749 140
rect 751 138 759 140
rect 747 134 759 138
rect 779 147 783 156
rect 770 146 783 147
rect 770 144 775 146
rect 777 144 783 146
rect 770 142 783 144
rect 892 129 902 216
rect 71 128 902 129
rect 931 128 939 129
rect 71 126 167 128
rect 169 126 195 128
rect 197 126 391 128
rect 393 126 419 128
rect 421 126 615 128
rect 617 126 643 128
rect 645 126 750 128
rect 752 126 760 128
rect 762 126 939 128
rect 71 121 939 126
rect 232 120 238 121
rect 780 120 901 121
rect 780 119 896 120
rect 29 94 913 99
rect 29 92 77 94
rect 79 92 91 94
rect 93 92 105 94
rect 107 92 210 94
rect 212 92 344 94
rect 346 92 358 94
rect 360 92 372 94
rect 374 92 476 94
rect 478 92 611 94
rect 613 92 625 94
rect 627 92 639 94
rect 641 92 742 94
rect 744 92 876 94
rect 878 92 890 94
rect 892 92 904 94
rect 906 92 913 94
rect 29 91 913 92
rect 74 69 78 78
rect 74 67 76 69
rect 74 46 78 67
rect 89 84 102 86
rect 89 82 93 84
rect 95 82 102 84
rect 89 80 102 82
rect 89 73 95 80
rect 118 81 131 85
rect 207 82 220 85
rect 118 79 123 81
rect 118 77 120 79
rect 122 77 123 79
rect 207 80 209 82
rect 211 81 220 82
rect 247 81 260 85
rect 118 72 123 77
rect 118 70 120 72
rect 122 70 123 72
rect 118 68 123 70
rect 74 44 76 46
rect 78 44 86 46
rect 74 40 86 44
rect 106 53 110 62
rect 97 52 110 53
rect 97 50 102 52
rect 104 50 110 52
rect 97 48 110 50
rect 118 46 122 68
rect 149 65 187 69
rect 149 62 154 65
rect 146 60 154 62
rect 146 58 147 60
rect 149 58 154 60
rect 146 56 154 58
rect 164 60 179 61
rect 164 58 166 60
rect 168 58 173 60
rect 175 58 179 60
rect 164 57 179 58
rect 118 44 123 46
rect 166 51 170 57
rect 197 76 203 78
rect 197 74 198 76
rect 200 74 203 76
rect 197 69 203 74
rect 197 67 198 69
rect 200 67 203 69
rect 197 65 203 67
rect 166 49 167 51
rect 169 49 170 51
rect 166 48 170 49
rect 199 45 203 65
rect 118 42 120 44
rect 122 42 123 44
rect 118 40 123 42
rect 181 44 203 45
rect 181 42 198 44
rect 200 42 203 44
rect 181 41 203 42
rect 207 48 211 80
rect 247 79 252 81
rect 231 69 235 78
rect 247 77 249 79
rect 251 77 252 79
rect 247 72 252 77
rect 247 70 249 72
rect 251 70 252 72
rect 222 68 235 69
rect 222 66 223 68
rect 225 66 226 68
rect 228 66 235 68
rect 222 65 235 66
rect 239 69 243 70
rect 239 67 240 69
rect 242 67 243 69
rect 239 61 243 67
rect 230 60 243 61
rect 230 58 236 60
rect 238 58 243 60
rect 230 57 243 58
rect 239 56 243 57
rect 247 68 252 70
rect 247 60 251 68
rect 247 58 248 60
rect 250 58 251 60
rect 278 65 316 69
rect 207 46 212 48
rect 207 44 209 46
rect 211 44 212 46
rect 70 34 202 35
rect 70 32 77 34
rect 79 32 87 34
rect 89 32 202 34
rect 70 31 202 32
rect 70 29 198 31
rect 200 29 202 31
rect 70 27 202 29
rect 207 10 212 44
rect 247 46 251 58
rect 278 62 283 65
rect 275 60 283 62
rect 275 58 276 60
rect 278 58 283 60
rect 275 56 283 58
rect 293 60 308 61
rect 293 58 295 60
rect 297 58 302 60
rect 304 58 308 60
rect 293 57 308 58
rect 295 53 299 57
rect 326 76 332 78
rect 326 74 327 76
rect 329 74 332 76
rect 326 69 332 74
rect 326 67 327 69
rect 329 67 332 69
rect 326 65 332 67
rect 247 44 252 46
rect 295 51 296 53
rect 298 51 299 53
rect 295 48 299 51
rect 328 45 332 65
rect 247 42 249 44
rect 251 42 252 44
rect 247 40 252 42
rect 310 44 332 45
rect 310 42 327 44
rect 329 42 332 44
rect 310 41 332 42
rect 341 69 345 78
rect 341 67 343 69
rect 341 53 345 67
rect 356 84 369 86
rect 356 82 360 84
rect 362 82 369 84
rect 356 80 369 82
rect 356 73 362 80
rect 384 81 397 85
rect 473 82 486 85
rect 384 79 389 81
rect 384 77 386 79
rect 388 77 389 79
rect 473 80 475 82
rect 477 81 486 82
rect 513 81 526 85
rect 384 72 389 77
rect 384 70 386 72
rect 388 70 389 72
rect 384 68 389 70
rect 341 51 342 53
rect 344 51 345 53
rect 341 46 345 51
rect 341 44 343 46
rect 345 44 353 46
rect 341 40 353 44
rect 373 53 377 62
rect 364 52 377 53
rect 364 50 369 52
rect 371 50 377 52
rect 364 48 377 50
rect 384 46 388 68
rect 415 65 453 69
rect 415 62 420 65
rect 412 60 420 62
rect 412 58 413 60
rect 415 58 420 60
rect 412 56 420 58
rect 430 60 445 61
rect 430 58 432 60
rect 434 58 439 60
rect 441 58 445 60
rect 430 57 445 58
rect 384 44 389 46
rect 432 51 436 57
rect 463 76 469 78
rect 463 74 464 76
rect 466 74 469 76
rect 463 69 469 74
rect 463 67 464 69
rect 466 67 469 69
rect 463 65 469 67
rect 432 49 433 51
rect 435 49 436 51
rect 432 48 436 49
rect 465 45 469 65
rect 384 42 386 44
rect 388 42 389 44
rect 384 40 389 42
rect 447 44 469 45
rect 447 42 464 44
rect 466 42 469 44
rect 447 41 469 42
rect 473 48 477 80
rect 513 79 518 81
rect 497 69 501 78
rect 513 77 515 79
rect 517 77 518 79
rect 513 72 518 77
rect 513 70 515 72
rect 517 70 518 72
rect 488 68 501 69
rect 488 66 489 68
rect 491 66 492 68
rect 494 66 501 68
rect 488 65 501 66
rect 505 69 509 70
rect 505 67 506 69
rect 508 67 509 69
rect 505 61 509 67
rect 496 60 509 61
rect 496 58 502 60
rect 504 58 509 60
rect 496 57 509 58
rect 505 56 509 57
rect 513 68 518 70
rect 513 60 517 68
rect 513 58 514 60
rect 516 58 517 60
rect 544 65 582 69
rect 473 46 478 48
rect 473 44 475 46
rect 477 44 478 46
rect 473 40 478 44
rect 217 34 464 35
rect 217 32 238 34
rect 240 32 344 34
rect 346 32 354 34
rect 356 32 464 34
rect 217 31 464 32
rect 217 29 219 31
rect 221 29 461 31
rect 463 29 464 31
rect 217 27 464 29
rect 473 13 477 40
rect 513 46 517 58
rect 544 62 549 65
rect 541 60 549 62
rect 541 58 542 60
rect 544 58 549 60
rect 541 56 549 58
rect 559 60 574 61
rect 559 58 561 60
rect 563 58 568 60
rect 570 58 574 60
rect 559 57 574 58
rect 513 44 518 46
rect 561 52 565 57
rect 592 76 598 78
rect 592 74 593 76
rect 595 74 598 76
rect 592 69 598 74
rect 592 67 593 69
rect 595 67 598 69
rect 592 65 598 67
rect 561 50 562 52
rect 564 50 565 52
rect 561 48 565 50
rect 594 45 598 65
rect 513 42 515 44
rect 517 42 518 44
rect 513 40 518 42
rect 576 44 598 45
rect 576 42 593 44
rect 595 42 598 44
rect 576 41 598 42
rect 608 69 612 78
rect 608 67 610 69
rect 608 52 612 67
rect 623 84 636 86
rect 623 82 627 84
rect 629 82 636 84
rect 623 80 636 82
rect 623 73 629 80
rect 650 81 663 85
rect 739 82 752 85
rect 650 79 655 81
rect 650 77 652 79
rect 654 77 655 79
rect 739 80 741 82
rect 743 81 752 82
rect 779 81 792 85
rect 650 72 655 77
rect 650 70 652 72
rect 654 70 655 72
rect 650 68 655 70
rect 608 50 609 52
rect 611 50 612 52
rect 608 46 612 50
rect 608 44 610 46
rect 612 44 620 46
rect 608 40 620 44
rect 640 53 644 62
rect 631 52 644 53
rect 631 50 636 52
rect 638 50 644 52
rect 631 48 644 50
rect 650 46 654 68
rect 681 68 719 69
rect 681 66 708 68
rect 710 66 719 68
rect 681 65 719 66
rect 681 62 686 65
rect 678 60 686 62
rect 678 58 679 60
rect 681 58 686 60
rect 678 56 686 58
rect 696 60 711 61
rect 696 58 698 60
rect 700 58 705 60
rect 707 58 711 60
rect 696 57 711 58
rect 650 44 655 46
rect 698 51 702 57
rect 729 76 735 78
rect 729 74 730 76
rect 732 74 735 76
rect 729 69 735 74
rect 729 67 730 69
rect 732 67 735 69
rect 729 65 735 67
rect 698 49 699 51
rect 701 49 702 51
rect 698 48 702 49
rect 731 45 735 65
rect 650 42 652 44
rect 654 42 655 44
rect 650 40 655 42
rect 713 44 735 45
rect 713 42 730 44
rect 732 42 735 44
rect 713 41 735 42
rect 739 48 743 80
rect 779 79 784 81
rect 763 69 767 78
rect 779 77 781 79
rect 783 77 784 79
rect 779 72 784 77
rect 779 70 781 72
rect 783 70 784 72
rect 754 68 767 69
rect 754 66 755 68
rect 757 66 758 68
rect 760 66 767 68
rect 754 65 767 66
rect 771 69 775 70
rect 771 67 772 69
rect 774 67 775 69
rect 771 61 775 67
rect 762 60 775 61
rect 762 58 768 60
rect 770 58 775 60
rect 762 57 775 58
rect 771 56 775 57
rect 779 68 784 70
rect 779 60 783 68
rect 779 58 780 60
rect 782 58 783 60
rect 810 65 848 69
rect 739 46 744 48
rect 739 44 741 46
rect 743 44 744 46
rect 739 41 744 44
rect 482 34 732 35
rect 482 32 504 34
rect 506 32 611 34
rect 613 32 621 34
rect 623 32 732 34
rect 482 31 732 32
rect 482 29 487 31
rect 489 29 729 31
rect 731 29 732 31
rect 482 27 732 29
rect 472 12 477 13
rect 739 16 743 41
rect 779 46 783 58
rect 810 62 815 65
rect 807 60 815 62
rect 807 58 808 60
rect 810 58 815 60
rect 807 56 815 58
rect 825 60 840 61
rect 825 58 827 60
rect 829 58 834 60
rect 836 58 840 60
rect 825 57 840 58
rect 779 44 784 46
rect 827 51 831 57
rect 858 76 864 78
rect 858 74 859 76
rect 861 74 864 76
rect 858 69 864 74
rect 858 67 859 69
rect 861 67 864 69
rect 858 65 864 67
rect 827 49 828 51
rect 830 49 831 51
rect 827 48 831 49
rect 860 45 864 65
rect 779 42 781 44
rect 783 42 784 44
rect 779 40 784 42
rect 842 44 864 45
rect 842 42 859 44
rect 861 42 864 44
rect 842 41 864 42
rect 873 69 877 78
rect 873 67 875 69
rect 873 52 877 67
rect 888 84 901 86
rect 888 82 892 84
rect 894 82 901 84
rect 888 80 901 82
rect 888 73 894 80
rect 873 50 874 52
rect 876 50 877 52
rect 873 46 877 50
rect 873 44 875 46
rect 877 44 885 46
rect 873 40 885 44
rect 905 53 909 62
rect 896 52 909 53
rect 896 50 901 52
rect 903 50 909 52
rect 896 48 909 50
rect 748 34 913 35
rect 931 34 939 121
rect 748 32 770 34
rect 772 32 876 34
rect 878 32 886 34
rect 888 32 939 34
rect 748 30 757 32
rect 759 30 939 32
rect 748 28 939 30
rect 748 27 913 28
rect 931 27 939 28
rect 739 14 740 16
rect 742 14 743 16
rect 739 12 743 14
rect 472 10 473 12
rect 475 10 477 12
rect 472 8 477 10
<< alu2 >>
rect 174 423 583 424
rect 883 423 894 424
rect 174 415 894 423
rect 174 414 583 415
rect 174 366 182 414
rect 867 404 876 405
rect 404 397 876 404
rect 174 364 176 366
rect 178 364 182 366
rect 174 363 182 364
rect 231 386 398 391
rect 231 350 237 386
rect 231 348 234 350
rect 236 348 237 350
rect 231 347 237 348
rect 254 351 260 352
rect 296 351 387 352
rect 254 349 255 351
rect 257 350 283 351
rect 257 349 280 350
rect 254 348 280 349
rect 282 348 283 350
rect 296 349 297 351
rect 299 349 384 351
rect 386 349 387 351
rect 296 348 387 349
rect 254 347 283 348
rect 54 343 80 344
rect 167 343 172 344
rect 392 343 398 386
rect 404 366 412 397
rect 404 364 407 366
rect 409 364 412 366
rect 404 363 412 364
rect 456 382 708 389
rect 456 350 461 382
rect 703 354 708 382
rect 741 384 746 386
rect 741 382 743 384
rect 745 382 746 384
rect 741 366 746 382
rect 741 364 742 366
rect 744 364 746 366
rect 741 363 746 364
rect 790 384 795 386
rect 790 382 792 384
rect 794 382 795 384
rect 790 366 795 382
rect 790 364 791 366
rect 793 364 795 366
rect 790 362 795 364
rect 840 384 845 386
rect 840 382 842 384
rect 844 382 845 384
rect 840 366 845 382
rect 840 364 841 366
rect 843 364 845 366
rect 840 362 845 364
rect 703 352 705 354
rect 707 352 708 354
rect 456 348 458 350
rect 460 348 461 350
rect 456 347 461 348
rect 478 351 484 352
rect 520 351 611 352
rect 478 349 479 351
rect 481 350 507 351
rect 481 349 504 350
rect 478 348 504 349
rect 506 348 507 350
rect 520 349 521 351
rect 523 349 608 351
rect 610 349 611 351
rect 520 348 611 349
rect 703 348 708 352
rect 478 347 507 348
rect 54 341 76 343
rect 78 341 80 343
rect 54 339 80 341
rect 103 342 108 343
rect 103 340 104 342
rect 106 340 108 342
rect 54 202 62 339
rect 103 306 108 340
rect 167 342 268 343
rect 167 340 265 342
rect 267 340 268 342
rect 167 339 268 340
rect 300 342 309 343
rect 300 340 305 342
rect 307 340 309 342
rect 300 339 309 340
rect 332 342 337 343
rect 332 340 333 342
rect 335 340 337 342
rect 167 335 172 339
rect 156 334 172 335
rect 123 333 172 334
rect 123 331 124 333
rect 126 331 172 333
rect 223 333 266 334
rect 300 333 304 339
rect 223 331 224 333
rect 226 331 304 333
rect 123 330 160 331
rect 223 330 304 331
rect 262 328 304 330
rect 138 325 166 326
rect 138 323 162 325
rect 164 323 166 325
rect 138 322 166 323
rect 70 302 108 306
rect 154 304 161 322
rect 153 303 275 304
rect 70 246 74 302
rect 153 301 271 303
rect 273 301 275 303
rect 153 300 275 301
rect 153 299 259 300
rect 268 299 275 300
rect 332 297 337 340
rect 392 342 492 343
rect 392 340 489 342
rect 491 340 492 342
rect 392 339 492 340
rect 524 342 533 343
rect 524 340 529 342
rect 531 340 533 342
rect 524 339 533 340
rect 556 342 564 343
rect 556 340 561 342
rect 563 340 564 342
rect 392 338 488 339
rect 319 293 337 297
rect 352 334 356 335
rect 352 332 353 334
rect 355 332 356 334
rect 352 297 356 332
rect 447 333 490 334
rect 524 333 528 339
rect 556 338 564 340
rect 652 341 659 342
rect 652 339 656 341
rect 658 339 659 341
rect 447 331 448 333
rect 450 331 528 333
rect 447 330 528 331
rect 486 328 528 330
rect 557 300 561 338
rect 352 293 372 297
rect 92 290 98 291
rect 92 288 94 290
rect 96 288 98 290
rect 92 272 98 288
rect 92 270 94 272
rect 96 270 98 272
rect 92 268 98 270
rect 142 290 148 291
rect 142 288 144 290
rect 146 288 148 290
rect 142 272 148 288
rect 142 270 144 272
rect 146 270 148 272
rect 142 268 148 270
rect 119 247 129 249
rect 70 245 79 246
rect 70 243 76 245
rect 78 243 79 245
rect 119 245 121 247
rect 123 245 126 247
rect 128 245 129 247
rect 119 244 129 245
rect 319 246 324 293
rect 342 277 348 279
rect 342 275 344 277
rect 346 275 348 277
rect 342 272 348 275
rect 342 270 344 272
rect 346 270 348 272
rect 342 268 348 270
rect 368 248 372 293
rect 519 296 561 300
rect 576 333 580 334
rect 576 331 577 333
rect 579 331 580 333
rect 576 296 580 331
rect 652 300 659 339
rect 772 338 776 341
rect 672 336 727 337
rect 672 335 724 336
rect 672 333 673 335
rect 675 334 724 335
rect 726 334 727 336
rect 675 333 727 334
rect 672 332 727 333
rect 772 336 773 338
rect 775 336 776 338
rect 437 291 443 292
rect 437 289 439 291
rect 441 289 443 291
rect 437 288 443 289
rect 392 272 403 274
rect 392 270 394 272
rect 396 270 400 272
rect 402 270 403 272
rect 392 268 403 270
rect 437 272 441 288
rect 437 270 438 272
rect 440 270 441 272
rect 437 269 441 270
rect 492 272 515 274
rect 492 270 494 272
rect 496 270 500 272
rect 502 270 512 272
rect 514 270 515 272
rect 492 268 515 270
rect 368 247 379 248
rect 319 244 329 246
rect 368 245 376 247
rect 378 245 379 247
rect 368 244 379 245
rect 519 244 524 296
rect 571 292 580 296
rect 621 296 659 300
rect 772 296 776 336
rect 822 337 826 342
rect 822 335 823 337
rect 825 335 826 337
rect 822 296 826 335
rect 528 272 548 274
rect 528 270 529 272
rect 531 270 544 272
rect 546 270 548 272
rect 528 268 548 270
rect 571 245 575 292
rect 591 272 603 274
rect 591 270 594 272
rect 596 270 600 272
rect 602 270 603 272
rect 591 268 603 270
rect 621 247 625 296
rect 700 292 776 296
rect 800 292 826 296
rect 629 272 654 274
rect 629 270 630 272
rect 632 270 650 272
rect 652 270 654 272
rect 629 268 654 270
rect 700 248 704 292
rect 621 246 629 247
rect 571 244 579 245
rect 70 242 79 243
rect 319 242 326 244
rect 328 242 329 244
rect 519 243 529 244
rect 319 241 329 242
rect 475 241 479 243
rect 475 239 476 241
rect 478 239 479 241
rect 519 241 526 243
rect 528 241 529 243
rect 571 242 576 244
rect 578 242 579 244
rect 621 244 626 246
rect 628 244 629 246
rect 700 246 701 248
rect 703 246 704 248
rect 700 245 704 246
rect 716 248 722 249
rect 716 246 717 248
rect 719 246 722 248
rect 621 243 629 244
rect 571 241 579 242
rect 519 240 529 241
rect 53 120 62 202
rect 75 209 80 211
rect 75 207 76 209
rect 78 207 80 209
rect 75 157 80 207
rect 131 209 396 213
rect 475 212 479 239
rect 475 210 476 212
rect 478 210 479 212
rect 475 209 479 210
rect 716 212 722 246
rect 800 248 804 292
rect 800 246 801 248
rect 803 246 804 248
rect 800 245 804 246
rect 816 239 821 248
rect 816 237 818 239
rect 820 237 821 239
rect 716 210 718 212
rect 720 210 722 212
rect 131 205 140 209
rect 131 159 139 205
rect 387 203 396 209
rect 612 208 618 209
rect 497 204 618 208
rect 716 207 722 210
rect 748 232 754 235
rect 748 230 749 232
rect 751 230 754 232
rect 748 212 754 230
rect 748 210 750 212
rect 752 210 754 212
rect 748 209 754 210
rect 816 205 821 237
rect 284 201 295 202
rect 284 199 291 201
rect 293 199 295 201
rect 284 198 295 199
rect 164 197 168 198
rect 164 195 165 197
rect 167 195 168 197
rect 164 179 168 195
rect 164 175 175 179
rect 164 171 168 175
rect 164 169 165 171
rect 167 169 168 171
rect 164 168 168 169
rect 154 163 160 164
rect 196 163 287 164
rect 154 161 155 163
rect 157 162 183 163
rect 157 161 180 162
rect 154 160 180 161
rect 182 160 183 162
rect 196 161 197 163
rect 199 161 284 163
rect 286 161 287 163
rect 196 160 287 161
rect 154 159 183 160
rect 75 155 76 157
rect 78 155 80 157
rect 75 150 80 155
rect 200 154 209 155
rect 200 152 205 154
rect 207 152 209 154
rect 200 151 209 152
rect 232 154 238 155
rect 232 152 233 154
rect 235 152 238 154
rect 123 145 166 146
rect 200 145 204 151
rect 123 143 124 145
rect 126 143 204 145
rect 123 142 204 143
rect 162 140 204 142
rect 232 132 238 152
rect 291 149 295 198
rect 355 197 363 199
rect 355 195 358 197
rect 360 195 363 197
rect 355 159 363 195
rect 387 174 395 203
rect 497 198 504 204
rect 580 198 590 200
rect 439 197 504 198
rect 439 195 441 197
rect 443 195 504 197
rect 439 194 504 195
rect 516 197 520 198
rect 516 195 517 197
rect 519 195 520 197
rect 378 163 384 164
rect 420 163 511 164
rect 378 161 379 163
rect 381 162 407 163
rect 381 161 404 162
rect 378 160 404 161
rect 406 160 407 162
rect 420 161 421 163
rect 423 161 508 163
rect 510 161 511 163
rect 420 160 511 161
rect 378 159 407 160
rect 252 148 295 149
rect 252 146 253 148
rect 255 146 295 148
rect 424 154 433 155
rect 424 152 429 154
rect 431 152 433 154
rect 424 151 433 152
rect 456 154 460 155
rect 456 152 457 154
rect 459 152 460 154
rect 252 145 295 146
rect 232 130 234 132
rect 236 130 238 132
rect 232 128 238 130
rect 299 143 304 146
rect 299 141 300 143
rect 302 141 304 143
rect 347 145 390 146
rect 424 145 428 151
rect 347 143 348 145
rect 350 143 428 145
rect 347 142 428 143
rect 299 127 304 141
rect 386 140 428 142
rect 53 114 238 120
rect 298 119 304 127
rect 456 119 460 152
rect 516 149 520 195
rect 580 196 582 198
rect 584 196 590 198
rect 580 159 585 196
rect 612 172 618 204
rect 799 200 804 204
rect 816 203 817 205
rect 819 203 821 205
rect 816 201 821 203
rect 637 199 804 200
rect 637 197 639 199
rect 641 197 804 199
rect 637 196 804 197
rect 799 192 804 196
rect 849 192 854 265
rect 867 215 876 397
rect 868 205 876 215
rect 868 203 871 205
rect 873 203 876 205
rect 868 200 876 203
rect 799 188 854 192
rect 849 186 854 188
rect 883 192 894 415
rect 765 178 834 180
rect 765 176 766 178
rect 768 176 830 178
rect 832 176 834 178
rect 765 175 834 176
rect 602 163 608 164
rect 644 163 735 164
rect 602 161 603 163
rect 605 162 631 163
rect 605 161 628 162
rect 602 160 628 161
rect 630 160 631 162
rect 644 161 645 163
rect 647 161 732 163
rect 734 161 735 163
rect 644 160 735 161
rect 602 159 631 160
rect 476 148 520 149
rect 648 154 657 155
rect 648 152 653 154
rect 655 152 657 154
rect 648 151 657 152
rect 679 154 684 155
rect 679 152 681 154
rect 683 152 684 154
rect 476 146 477 148
rect 479 146 520 148
rect 476 144 520 146
rect 298 117 300 119
rect 302 117 304 119
rect 298 115 304 117
rect 232 110 238 114
rect 455 110 460 119
rect 232 105 460 110
rect 524 138 529 148
rect 571 145 614 146
rect 648 145 652 151
rect 571 143 572 145
rect 574 143 652 145
rect 571 142 652 143
rect 610 140 652 142
rect 524 136 525 138
rect 527 136 529 138
rect 524 104 529 136
rect 679 118 684 152
rect 699 146 751 148
rect 699 144 701 146
rect 703 144 748 146
rect 750 144 751 146
rect 699 142 751 144
rect 883 118 892 192
rect 678 113 898 118
rect 883 112 892 113
rect 524 102 525 104
rect 527 102 529 104
rect 524 101 529 102
rect 625 86 631 111
rect 707 102 796 104
rect 707 100 790 102
rect 792 100 796 102
rect 707 99 796 100
rect 891 103 896 104
rect 891 101 893 103
rect 895 101 896 103
rect 343 84 364 86
rect 343 82 345 84
rect 347 82 360 84
rect 362 82 364 84
rect 343 80 364 82
rect 608 84 631 86
rect 608 82 610 84
rect 612 82 627 84
rect 629 82 631 84
rect 608 80 631 82
rect 197 69 203 70
rect 239 69 330 70
rect 197 67 198 69
rect 200 68 226 69
rect 200 67 223 68
rect 197 66 223 67
rect 225 66 226 68
rect 239 67 240 69
rect 242 67 327 69
rect 329 67 330 69
rect 239 66 330 67
rect 463 69 469 70
rect 505 69 596 70
rect 463 67 464 69
rect 466 68 492 69
rect 466 67 489 68
rect 463 66 489 67
rect 491 66 492 68
rect 505 67 506 69
rect 508 67 593 69
rect 595 67 596 69
rect 505 66 596 67
rect 706 68 712 99
rect 891 84 896 101
rect 891 82 892 84
rect 894 82 896 84
rect 891 80 896 82
rect 706 66 708 68
rect 710 66 712 68
rect 197 65 226 66
rect 463 65 492 66
rect 706 65 712 66
rect 729 69 735 70
rect 771 69 862 70
rect 729 67 730 69
rect 732 68 758 69
rect 732 67 755 68
rect 729 66 755 67
rect 757 66 758 68
rect 771 67 772 69
rect 774 67 859 69
rect 861 67 862 69
rect 771 66 862 67
rect 729 65 758 66
rect 146 60 151 62
rect 146 58 147 60
rect 149 58 151 60
rect 146 8 151 58
rect 243 60 252 61
rect 243 58 248 60
rect 250 58 252 60
rect 243 57 252 58
rect 274 60 281 62
rect 274 58 276 60
rect 278 58 281 60
rect 166 51 209 52
rect 243 51 247 57
rect 166 49 167 51
rect 169 49 247 51
rect 166 48 247 49
rect 205 46 247 48
rect 196 31 224 34
rect 196 29 198 31
rect 200 29 219 31
rect 221 29 224 31
rect 196 27 224 29
rect 274 22 281 58
rect 412 60 418 62
rect 412 58 413 60
rect 415 58 418 60
rect 295 53 345 55
rect 295 51 296 53
rect 298 51 342 53
rect 344 51 345 53
rect 295 50 345 51
rect 274 20 277 22
rect 279 20 281 22
rect 274 19 281 20
rect 145 -4 151 8
rect 145 -6 146 -4
rect 148 -6 151 -4
rect 145 -8 151 -6
rect 412 0 418 58
rect 509 60 518 61
rect 509 58 514 60
rect 516 58 518 60
rect 509 57 518 58
rect 541 60 547 62
rect 541 58 542 60
rect 544 58 547 60
rect 432 51 475 52
rect 509 51 513 57
rect 432 49 433 51
rect 435 49 513 51
rect 432 48 513 49
rect 471 46 513 48
rect 458 31 492 35
rect 458 29 461 31
rect 463 29 487 31
rect 489 29 492 31
rect 458 27 492 29
rect 541 26 547 58
rect 775 60 784 61
rect 775 58 780 60
rect 782 58 784 60
rect 775 57 784 58
rect 807 60 812 62
rect 807 58 808 60
rect 810 58 812 60
rect 561 52 612 53
rect 561 50 562 52
rect 564 50 609 52
rect 611 50 612 52
rect 561 48 612 50
rect 698 51 741 52
rect 775 51 779 57
rect 698 49 699 51
rect 701 49 779 51
rect 698 48 779 49
rect 737 46 779 48
rect 726 32 761 35
rect 726 31 757 32
rect 726 29 729 31
rect 731 30 757 31
rect 759 30 761 32
rect 731 29 761 30
rect 726 27 761 29
rect 540 20 548 26
rect 540 18 543 20
rect 545 18 548 20
rect 540 17 548 18
rect 448 12 477 14
rect 448 10 450 12
rect 452 10 473 12
rect 475 10 477 12
rect 448 8 477 10
rect 497 13 637 17
rect 497 11 500 13
rect 502 12 637 13
rect 502 11 631 12
rect 497 10 631 11
rect 633 10 637 12
rect 497 7 637 10
rect 738 16 743 17
rect 738 14 740 16
rect 742 14 743 16
rect 738 0 743 14
rect 412 -7 746 0
rect 807 -18 812 58
rect 827 52 877 53
rect 827 51 874 52
rect 827 49 828 51
rect 830 50 874 51
rect 876 50 877 52
rect 830 49 877 50
rect 827 48 877 49
rect 807 -20 808 -18
rect 810 -20 812 -18
rect 807 -22 812 -20
<< alu3 >>
rect 436 425 847 431
rect 92 384 348 387
rect 92 382 335 384
rect 337 382 348 384
rect 92 381 348 382
rect 92 290 98 381
rect 92 288 94 290
rect 96 288 98 290
rect 92 286 98 288
rect 142 290 148 381
rect 142 288 144 290
rect 146 288 148 290
rect 142 287 148 288
rect 268 303 277 304
rect 268 301 271 303
rect 273 301 277 303
rect 120 247 124 249
rect 120 245 121 247
rect 123 245 124 247
rect 120 232 124 245
rect 120 228 208 232
rect 37 209 80 211
rect 37 207 76 209
rect 78 207 80 209
rect 37 206 80 207
rect 37 17 41 206
rect 54 197 168 198
rect 54 195 165 197
rect 167 195 168 197
rect 54 193 168 195
rect 54 23 65 193
rect 204 134 208 228
rect 268 203 277 301
rect 342 277 348 381
rect 437 291 443 425
rect 741 384 747 425
rect 741 382 743 384
rect 745 382 747 384
rect 741 381 747 382
rect 790 384 795 425
rect 790 382 792 384
rect 794 382 795 384
rect 840 384 846 425
rect 840 382 842 384
rect 844 382 846 384
rect 790 381 795 382
rect 841 381 846 382
rect 437 289 439 291
rect 441 289 443 291
rect 437 288 443 289
rect 342 275 344 277
rect 346 275 348 277
rect 342 274 348 275
rect 398 272 532 274
rect 398 270 400 272
rect 402 270 500 272
rect 502 270 512 272
rect 514 270 529 272
rect 531 270 532 272
rect 398 268 532 270
rect 598 272 917 274
rect 598 270 600 272
rect 602 270 630 272
rect 632 270 917 272
rect 598 268 917 270
rect 475 212 479 215
rect 475 210 476 212
rect 478 210 479 212
rect 267 201 296 203
rect 267 199 291 201
rect 293 199 296 201
rect 267 196 296 199
rect 475 198 479 210
rect 510 213 516 268
rect 618 267 917 268
rect 510 212 604 213
rect 510 210 601 212
rect 603 210 604 212
rect 510 208 604 210
rect 716 212 723 214
rect 716 210 718 212
rect 720 210 723 212
rect 580 199 648 200
rect 580 198 639 199
rect 355 197 445 198
rect 355 195 358 197
rect 360 195 441 197
rect 443 195 445 197
rect 355 194 445 195
rect 475 197 520 198
rect 475 195 517 197
rect 519 195 520 197
rect 580 196 582 198
rect 584 197 639 198
rect 641 197 648 199
rect 584 196 648 197
rect 580 195 648 196
rect 475 194 520 195
rect 233 134 238 135
rect 204 132 238 134
rect 204 130 234 132
rect 236 130 238 132
rect 204 129 238 130
rect 298 119 304 126
rect 298 117 300 119
rect 302 117 304 119
rect 298 104 304 117
rect 716 106 723 210
rect 748 212 754 214
rect 748 210 750 212
rect 752 210 795 212
rect 748 208 795 210
rect 497 104 505 106
rect 298 99 505 104
rect 524 104 723 106
rect 524 102 525 104
rect 527 102 723 104
rect 524 100 723 102
rect 716 99 723 100
rect 788 110 795 208
rect 815 205 876 208
rect 815 203 817 205
rect 819 203 871 205
rect 873 203 876 205
rect 815 201 876 203
rect 827 178 834 180
rect 827 176 830 178
rect 832 176 834 178
rect 788 102 796 110
rect 788 100 790 102
rect 792 100 796 102
rect 827 104 834 176
rect 908 105 917 267
rect 884 104 918 105
rect 827 103 918 104
rect 827 101 893 103
rect 895 101 918 103
rect 827 100 918 101
rect 788 99 796 100
rect 884 99 918 100
rect 334 84 356 86
rect 334 82 337 84
rect 339 82 345 84
rect 347 82 356 84
rect 334 80 356 82
rect 54 22 282 23
rect 54 20 277 22
rect 279 20 282 22
rect 36 -23 42 17
rect 54 16 282 20
rect 348 12 455 14
rect 348 10 450 12
rect 452 10 455 12
rect 348 8 455 10
rect 497 13 505 99
rect 599 84 614 86
rect 599 82 601 84
rect 603 82 610 84
rect 612 82 614 84
rect 599 80 614 82
rect 747 37 755 99
rect 497 11 500 13
rect 502 11 505 13
rect 497 8 505 11
rect 540 20 548 26
rect 748 23 755 37
rect 540 18 543 20
rect 545 18 548 20
rect 348 0 356 8
rect 145 -4 356 0
rect 145 -6 146 -4
rect 148 -6 356 -4
rect 145 -8 356 -6
rect 348 -9 356 -8
rect 540 -23 548 18
rect 629 12 636 17
rect 629 10 631 12
rect 633 10 636 12
rect 629 -16 636 10
rect 628 -18 812 -16
rect 628 -20 808 -18
rect 810 -20 812 -18
rect 628 -22 812 -20
rect 36 -32 548 -23
rect 36 -33 42 -32
<< alu4 >>
rect 333 384 340 395
rect 333 382 335 384
rect 337 382 340 384
rect 333 86 340 382
rect 599 212 604 213
rect 599 210 601 212
rect 603 210 604 212
rect 331 84 345 86
rect 331 82 337 84
rect 339 82 345 84
rect 331 80 345 82
rect 599 84 604 210
rect 599 82 601 84
rect 603 82 604 84
rect 599 80 604 82
<< ptie >>
rect 265 316 299 318
rect 265 314 267 316
rect 269 314 295 316
rect 297 314 299 316
rect 265 312 299 314
rect 489 316 523 318
rect 489 314 491 316
rect 493 314 519 316
rect 521 314 523 316
rect 489 312 523 314
rect 724 316 730 318
rect 724 314 726 316
rect 728 314 730 316
rect 724 312 730 314
rect 773 316 779 318
rect 773 314 775 316
rect 777 314 779 316
rect 773 312 779 314
rect 823 316 829 318
rect 823 314 825 316
rect 827 314 829 316
rect 823 312 829 314
rect 76 222 82 224
rect 76 220 78 222
rect 80 220 82 222
rect 76 218 82 220
rect 126 222 132 224
rect 126 220 128 222
rect 130 220 132 222
rect 126 218 132 220
rect 197 223 203 225
rect 197 221 199 223
rect 201 221 203 223
rect 197 219 203 221
rect 238 223 244 225
rect 238 221 240 223
rect 242 221 244 223
rect 238 219 244 221
rect 326 222 332 224
rect 326 220 328 222
rect 330 220 332 222
rect 326 218 332 220
rect 376 222 382 224
rect 376 220 378 222
rect 380 220 382 222
rect 376 218 382 220
rect 420 222 426 224
rect 420 220 422 222
rect 424 220 426 222
rect 420 218 426 220
rect 476 222 482 224
rect 476 220 478 222
rect 480 220 482 222
rect 476 218 482 220
rect 526 222 532 224
rect 526 220 528 222
rect 530 220 532 222
rect 526 218 532 220
rect 576 222 582 224
rect 576 220 578 222
rect 580 220 582 222
rect 576 218 582 220
rect 626 222 632 224
rect 626 220 628 222
rect 630 220 632 222
rect 626 218 632 220
rect 165 128 199 130
rect 165 126 167 128
rect 169 126 195 128
rect 197 126 199 128
rect 165 124 199 126
rect 389 128 423 130
rect 389 126 391 128
rect 393 126 419 128
rect 421 126 423 128
rect 389 124 423 126
rect 613 128 647 130
rect 613 126 615 128
rect 617 126 643 128
rect 645 126 647 128
rect 613 124 647 126
rect 748 128 754 130
rect 748 126 750 128
rect 752 126 754 128
rect 748 124 754 126
rect 75 34 81 36
rect 75 32 77 34
rect 79 32 81 34
rect 75 30 81 32
rect 217 34 242 36
rect 217 32 238 34
rect 240 32 242 34
rect 217 30 242 32
rect 342 34 348 36
rect 342 32 344 34
rect 346 32 348 34
rect 342 30 348 32
rect 482 34 508 36
rect 482 32 504 34
rect 506 32 508 34
rect 482 30 508 32
rect 609 34 615 36
rect 609 32 611 34
rect 613 32 615 34
rect 609 30 615 32
rect 748 34 774 36
rect 748 32 770 34
rect 772 32 774 34
rect 748 30 774 32
rect 874 34 880 36
rect 874 32 876 34
rect 878 32 880 34
rect 874 30 880 32
<< ntie >>
rect 265 376 271 378
rect 265 374 267 376
rect 269 374 271 376
rect 265 372 271 374
rect 489 376 495 378
rect 489 374 491 376
rect 493 374 495 376
rect 489 372 495 374
rect 724 376 758 378
rect 724 374 726 376
rect 728 374 740 376
rect 742 374 754 376
rect 756 374 758 376
rect 724 372 758 374
rect 773 376 807 378
rect 773 374 775 376
rect 777 374 789 376
rect 791 374 803 376
rect 805 374 807 376
rect 773 372 807 374
rect 823 376 857 378
rect 823 374 825 376
rect 827 374 839 376
rect 841 374 853 376
rect 855 374 857 376
rect 823 372 857 374
rect 76 282 110 284
rect 76 280 78 282
rect 80 280 92 282
rect 94 280 106 282
rect 108 280 110 282
rect 76 278 110 280
rect 126 282 160 284
rect 126 280 128 282
rect 130 280 142 282
rect 144 280 156 282
rect 158 280 160 282
rect 126 278 160 280
rect 197 283 231 285
rect 197 281 199 283
rect 201 281 213 283
rect 215 281 227 283
rect 229 281 231 283
rect 197 279 231 281
rect 238 283 272 285
rect 238 281 240 283
rect 242 281 254 283
rect 256 281 268 283
rect 270 281 272 283
rect 238 279 272 281
rect 326 282 360 284
rect 326 280 328 282
rect 330 280 342 282
rect 344 280 356 282
rect 358 280 360 282
rect 326 278 360 280
rect 376 282 410 284
rect 376 280 378 282
rect 380 280 392 282
rect 394 280 406 282
rect 408 280 410 282
rect 376 278 410 280
rect 420 282 454 284
rect 420 280 422 282
rect 424 280 436 282
rect 438 280 450 282
rect 452 280 454 282
rect 420 278 454 280
rect 476 282 510 284
rect 476 280 478 282
rect 480 280 492 282
rect 494 280 506 282
rect 508 280 510 282
rect 476 278 510 280
rect 526 282 560 284
rect 526 280 528 282
rect 530 280 542 282
rect 544 280 556 282
rect 558 280 560 282
rect 526 278 560 280
rect 576 282 610 284
rect 576 280 578 282
rect 580 280 592 282
rect 594 280 606 282
rect 608 280 610 282
rect 576 278 610 280
rect 626 282 660 284
rect 626 280 628 282
rect 630 280 642 282
rect 644 280 656 282
rect 658 280 660 282
rect 626 278 660 280
rect 165 188 171 190
rect 165 186 167 188
rect 169 186 171 188
rect 165 184 171 186
rect 389 188 395 190
rect 389 186 391 188
rect 393 186 395 188
rect 389 184 395 186
rect 613 188 619 190
rect 613 186 615 188
rect 617 186 619 188
rect 613 184 619 186
rect 748 188 782 190
rect 748 186 750 188
rect 752 186 764 188
rect 766 186 778 188
rect 780 186 782 188
rect 748 184 782 186
rect 75 94 109 96
rect 75 92 77 94
rect 79 92 91 94
rect 93 92 105 94
rect 107 92 109 94
rect 75 90 109 92
rect 208 94 214 96
rect 208 92 210 94
rect 212 92 214 94
rect 208 90 214 92
rect 342 94 376 96
rect 342 92 344 94
rect 346 92 358 94
rect 360 92 372 94
rect 374 92 376 94
rect 342 90 376 92
rect 474 94 480 96
rect 474 92 476 94
rect 478 92 480 94
rect 474 90 480 92
rect 609 94 643 96
rect 609 92 611 94
rect 613 92 625 94
rect 627 92 639 94
rect 641 92 643 94
rect 609 90 643 92
rect 740 94 746 96
rect 740 92 742 94
rect 744 92 746 94
rect 740 90 746 92
rect 874 94 908 96
rect 874 92 876 94
rect 878 92 890 94
rect 892 92 904 94
rect 906 92 908 94
rect 874 90 908 92
<< nmos >>
rect 82 315 84 328
rect 92 318 94 328
rect 102 321 104 335
rect 112 321 114 335
rect 132 315 134 335
rect 139 315 141 335
rect 150 315 152 329
rect 182 315 184 328
rect 192 318 194 328
rect 202 321 204 335
rect 212 321 214 335
rect 232 315 234 335
rect 239 315 241 335
rect 250 315 252 329
rect 271 324 273 330
rect 281 324 283 330
rect 291 324 293 330
rect 311 315 313 328
rect 321 318 323 328
rect 331 321 333 335
rect 341 321 343 335
rect 361 315 363 335
rect 368 315 370 335
rect 379 315 381 329
rect 406 315 408 328
rect 416 318 418 328
rect 426 321 428 335
rect 436 321 438 335
rect 456 315 458 335
rect 463 315 465 335
rect 474 315 476 329
rect 495 324 497 330
rect 505 324 507 330
rect 515 324 517 330
rect 535 315 537 328
rect 545 318 547 328
rect 555 321 557 335
rect 565 321 567 335
rect 585 315 587 335
rect 592 315 594 335
rect 603 315 605 329
rect 631 315 633 328
rect 641 318 643 328
rect 651 321 653 335
rect 661 321 663 335
rect 681 315 683 335
rect 688 315 690 335
rect 699 315 701 329
rect 730 324 732 330
rect 742 318 744 327
rect 749 318 751 327
rect 779 324 781 330
rect 791 318 793 327
rect 798 318 800 327
rect 829 324 831 330
rect 841 318 843 327
rect 848 318 850 327
rect 82 230 84 236
rect 94 224 96 233
rect 101 224 103 233
rect 132 230 134 236
rect 144 224 146 233
rect 151 224 153 233
rect 203 231 205 237
rect 215 225 217 234
rect 222 225 224 234
rect 244 231 246 237
rect 256 225 258 234
rect 263 225 265 234
rect 332 230 334 236
rect 344 224 346 233
rect 351 224 353 233
rect 382 230 384 236
rect 394 224 396 233
rect 401 224 403 233
rect 426 230 428 236
rect 438 224 440 233
rect 445 224 447 233
rect 482 230 484 236
rect 494 224 496 233
rect 501 224 503 233
rect 532 230 534 236
rect 544 224 546 233
rect 551 224 553 233
rect 582 230 584 236
rect 594 224 596 233
rect 601 224 603 233
rect 632 230 634 236
rect 644 224 646 233
rect 651 224 653 233
rect 676 221 678 234
rect 686 224 688 234
rect 696 227 698 241
rect 706 227 708 241
rect 726 221 728 241
rect 733 221 735 241
rect 744 221 746 235
rect 776 221 778 234
rect 786 224 788 234
rect 796 227 798 241
rect 806 227 808 241
rect 826 221 828 241
rect 833 221 835 241
rect 844 221 846 235
rect 82 127 84 140
rect 92 130 94 140
rect 102 133 104 147
rect 112 133 114 147
rect 132 127 134 147
rect 139 127 141 147
rect 150 127 152 141
rect 171 136 173 142
rect 181 136 183 142
rect 191 136 193 142
rect 211 127 213 140
rect 221 130 223 140
rect 231 133 233 147
rect 241 133 243 147
rect 261 127 263 147
rect 268 127 270 147
rect 279 127 281 141
rect 306 127 308 140
rect 316 130 318 140
rect 326 133 328 147
rect 336 133 338 147
rect 356 127 358 147
rect 363 127 365 147
rect 374 127 376 141
rect 395 136 397 142
rect 405 136 407 142
rect 415 136 417 142
rect 435 127 437 140
rect 445 130 447 140
rect 455 133 457 147
rect 465 133 467 147
rect 485 127 487 147
rect 492 127 494 147
rect 503 127 505 141
rect 530 127 532 140
rect 540 130 542 140
rect 550 133 552 147
rect 560 133 562 147
rect 580 127 582 147
rect 587 127 589 147
rect 598 127 600 141
rect 619 136 621 142
rect 629 136 631 142
rect 639 136 641 142
rect 659 127 661 140
rect 669 130 671 140
rect 679 133 681 147
rect 689 133 691 147
rect 709 127 711 147
rect 716 127 718 147
rect 727 127 729 141
rect 754 136 756 142
rect 766 130 768 139
rect 773 130 775 139
rect 81 42 83 48
rect 93 36 95 45
rect 100 36 102 45
rect 125 33 127 46
rect 135 36 137 46
rect 145 39 147 53
rect 155 39 157 53
rect 175 33 177 53
rect 182 33 184 53
rect 193 33 195 47
rect 214 42 216 48
rect 224 42 226 48
rect 234 42 236 48
rect 254 33 256 46
rect 264 36 266 46
rect 274 39 276 53
rect 284 39 286 53
rect 304 33 306 53
rect 311 33 313 53
rect 322 33 324 47
rect 348 42 350 48
rect 360 36 362 45
rect 367 36 369 45
rect 391 33 393 46
rect 401 36 403 46
rect 411 39 413 53
rect 421 39 423 53
rect 441 33 443 53
rect 448 33 450 53
rect 459 33 461 47
rect 480 42 482 48
rect 490 42 492 48
rect 500 42 502 48
rect 520 33 522 46
rect 530 36 532 46
rect 540 39 542 53
rect 550 39 552 53
rect 570 33 572 53
rect 577 33 579 53
rect 588 33 590 47
rect 615 42 617 48
rect 627 36 629 45
rect 634 36 636 45
rect 657 33 659 46
rect 667 36 669 46
rect 677 39 679 53
rect 687 39 689 53
rect 707 33 709 53
rect 714 33 716 53
rect 725 33 727 47
rect 746 42 748 48
rect 756 42 758 48
rect 766 42 768 48
rect 786 33 788 46
rect 796 36 798 46
rect 806 39 808 53
rect 816 39 818 53
rect 836 33 838 53
rect 843 33 845 53
rect 854 33 856 47
rect 880 42 882 48
rect 892 36 894 45
rect 899 36 901 45
<< pmos >>
rect 82 350 84 375
rect 95 350 97 363
rect 105 347 107 372
rect 112 347 114 372
rect 130 347 132 375
rect 140 347 142 375
rect 150 347 152 375
rect 182 350 184 375
rect 195 350 197 363
rect 205 347 207 372
rect 212 347 214 372
rect 230 347 232 375
rect 240 347 242 375
rect 250 347 252 375
rect 271 354 273 366
rect 284 357 286 375
rect 291 357 293 375
rect 311 350 313 375
rect 324 350 326 363
rect 334 347 336 372
rect 341 347 343 372
rect 359 347 361 375
rect 369 347 371 375
rect 379 347 381 375
rect 406 350 408 375
rect 419 350 421 363
rect 429 347 431 372
rect 436 347 438 372
rect 454 347 456 375
rect 464 347 466 375
rect 474 347 476 375
rect 495 354 497 366
rect 508 357 510 375
rect 515 357 517 375
rect 535 350 537 375
rect 548 350 550 363
rect 558 347 560 372
rect 565 347 567 372
rect 583 347 585 375
rect 593 347 595 375
rect 603 347 605 375
rect 631 350 633 375
rect 644 350 646 363
rect 654 347 656 372
rect 661 347 663 372
rect 679 347 681 375
rect 689 347 691 375
rect 699 347 701 375
rect 730 347 732 359
rect 740 347 742 357
rect 750 347 752 357
rect 779 347 781 359
rect 789 347 791 357
rect 799 347 801 357
rect 829 347 831 359
rect 839 347 841 357
rect 849 347 851 357
rect 82 253 84 265
rect 92 253 94 263
rect 102 253 104 263
rect 132 253 134 265
rect 142 253 144 263
rect 152 253 154 263
rect 203 254 205 266
rect 213 254 215 264
rect 223 254 225 264
rect 244 254 246 266
rect 254 254 256 264
rect 264 254 266 264
rect 332 253 334 265
rect 342 253 344 263
rect 352 253 354 263
rect 382 253 384 265
rect 392 253 394 263
rect 402 253 404 263
rect 426 253 428 265
rect 436 253 438 263
rect 446 253 448 263
rect 482 253 484 265
rect 492 253 494 263
rect 502 253 504 263
rect 532 253 534 265
rect 542 253 544 263
rect 552 253 554 263
rect 582 253 584 265
rect 592 253 594 263
rect 602 253 604 263
rect 632 253 634 265
rect 642 253 644 263
rect 652 253 654 263
rect 676 256 678 281
rect 689 256 691 269
rect 699 253 701 278
rect 706 253 708 278
rect 724 253 726 281
rect 734 253 736 281
rect 744 253 746 281
rect 776 256 778 281
rect 789 256 791 269
rect 799 253 801 278
rect 806 253 808 278
rect 824 253 826 281
rect 834 253 836 281
rect 844 253 846 281
rect 82 162 84 187
rect 95 162 97 175
rect 105 159 107 184
rect 112 159 114 184
rect 130 159 132 187
rect 140 159 142 187
rect 150 159 152 187
rect 171 166 173 178
rect 184 169 186 187
rect 191 169 193 187
rect 211 162 213 187
rect 224 162 226 175
rect 234 159 236 184
rect 241 159 243 184
rect 259 159 261 187
rect 269 159 271 187
rect 279 159 281 187
rect 306 162 308 187
rect 319 162 321 175
rect 329 159 331 184
rect 336 159 338 184
rect 354 159 356 187
rect 364 159 366 187
rect 374 159 376 187
rect 395 166 397 178
rect 408 169 410 187
rect 415 169 417 187
rect 435 162 437 187
rect 448 162 450 175
rect 458 159 460 184
rect 465 159 467 184
rect 483 159 485 187
rect 493 159 495 187
rect 503 159 505 187
rect 530 162 532 187
rect 543 162 545 175
rect 553 159 555 184
rect 560 159 562 184
rect 578 159 580 187
rect 588 159 590 187
rect 598 159 600 187
rect 619 166 621 178
rect 632 169 634 187
rect 639 169 641 187
rect 659 162 661 187
rect 672 162 674 175
rect 682 159 684 184
rect 689 159 691 184
rect 707 159 709 187
rect 717 159 719 187
rect 727 159 729 187
rect 754 159 756 171
rect 764 159 766 169
rect 774 159 776 169
rect 81 65 83 77
rect 91 65 93 75
rect 101 65 103 75
rect 125 68 127 93
rect 138 68 140 81
rect 148 65 150 90
rect 155 65 157 90
rect 173 65 175 93
rect 183 65 185 93
rect 193 65 195 93
rect 214 72 216 84
rect 227 75 229 93
rect 234 75 236 93
rect 254 68 256 93
rect 267 68 269 81
rect 277 65 279 90
rect 284 65 286 90
rect 302 65 304 93
rect 312 65 314 93
rect 322 65 324 93
rect 348 65 350 77
rect 358 65 360 75
rect 368 65 370 75
rect 391 68 393 93
rect 404 68 406 81
rect 414 65 416 90
rect 421 65 423 90
rect 439 65 441 93
rect 449 65 451 93
rect 459 65 461 93
rect 480 72 482 84
rect 493 75 495 93
rect 500 75 502 93
rect 520 68 522 93
rect 533 68 535 81
rect 543 65 545 90
rect 550 65 552 90
rect 568 65 570 93
rect 578 65 580 93
rect 588 65 590 93
rect 615 65 617 77
rect 625 65 627 75
rect 635 65 637 75
rect 657 68 659 93
rect 670 68 672 81
rect 680 65 682 90
rect 687 65 689 90
rect 705 65 707 93
rect 715 65 717 93
rect 725 65 727 93
rect 746 72 748 84
rect 759 75 761 93
rect 766 75 768 93
rect 786 68 788 93
rect 799 68 801 81
rect 809 65 811 90
rect 816 65 818 90
rect 834 65 836 93
rect 844 65 846 93
rect 854 65 856 93
rect 880 65 882 77
rect 890 65 892 75
rect 900 65 902 75
<< polyct0 >>
rect 90 343 92 345
rect 84 333 86 335
rect 140 340 142 342
rect 150 340 152 342
rect 190 343 192 345
rect 184 333 186 335
rect 240 340 242 342
rect 250 340 252 342
rect 273 341 275 343
rect 319 343 321 345
rect 313 333 315 335
rect 369 340 371 342
rect 379 340 381 342
rect 414 343 416 345
rect 408 333 410 335
rect 464 340 466 342
rect 474 340 476 342
rect 497 341 499 343
rect 543 343 545 345
rect 537 333 539 335
rect 593 340 595 342
rect 603 340 605 342
rect 639 343 641 345
rect 633 333 635 335
rect 689 340 691 342
rect 699 340 701 342
rect 732 340 734 342
rect 781 340 783 342
rect 831 340 833 342
rect 84 246 86 248
rect 134 246 136 248
rect 205 247 207 249
rect 246 247 248 249
rect 334 246 336 248
rect 384 246 386 248
rect 428 246 430 248
rect 484 246 486 248
rect 534 246 536 248
rect 584 246 586 248
rect 634 246 636 248
rect 684 249 686 251
rect 678 239 680 241
rect 734 246 736 248
rect 744 246 746 248
rect 784 249 786 251
rect 778 239 780 241
rect 834 246 836 248
rect 844 246 846 248
rect 90 155 92 157
rect 84 145 86 147
rect 140 152 142 154
rect 150 152 152 154
rect 173 153 175 155
rect 219 155 221 157
rect 213 145 215 147
rect 269 152 271 154
rect 279 152 281 154
rect 314 155 316 157
rect 308 145 310 147
rect 364 152 366 154
rect 374 152 376 154
rect 397 153 399 155
rect 443 155 445 157
rect 437 145 439 147
rect 493 152 495 154
rect 503 152 505 154
rect 538 155 540 157
rect 532 145 534 147
rect 588 152 590 154
rect 598 152 600 154
rect 621 153 623 155
rect 667 155 669 157
rect 661 145 663 147
rect 717 152 719 154
rect 727 152 729 154
rect 756 152 758 154
rect 83 58 85 60
rect 133 61 135 63
rect 127 51 129 53
rect 183 58 185 60
rect 193 58 195 60
rect 216 59 218 61
rect 262 61 264 63
rect 256 51 258 53
rect 312 58 314 60
rect 322 58 324 60
rect 350 58 352 60
rect 399 61 401 63
rect 393 51 395 53
rect 449 58 451 60
rect 459 58 461 60
rect 482 59 484 61
rect 528 61 530 63
rect 522 51 524 53
rect 578 58 580 60
rect 588 58 590 60
rect 617 58 619 60
rect 665 61 667 63
rect 659 51 661 53
rect 715 58 717 60
rect 725 58 727 60
rect 748 59 750 61
rect 794 61 796 63
rect 788 51 790 53
rect 844 58 846 60
rect 854 58 856 60
rect 882 58 884 60
<< polyct1 >>
rect 104 340 106 342
rect 123 340 125 342
rect 130 340 132 342
rect 283 348 285 350
rect 204 340 206 342
rect 223 340 225 342
rect 230 340 232 342
rect 293 340 295 342
rect 333 340 335 342
rect 352 340 354 342
rect 359 340 361 342
rect 507 348 509 350
rect 428 340 430 342
rect 447 340 449 342
rect 454 340 456 342
rect 517 340 519 342
rect 557 340 559 342
rect 576 340 578 342
rect 583 340 585 342
rect 742 364 744 366
rect 791 364 793 366
rect 841 364 843 366
rect 653 340 655 342
rect 672 340 674 342
rect 679 340 681 342
rect 751 332 753 334
rect 800 332 802 334
rect 850 332 852 334
rect 94 270 96 272
rect 144 270 146 272
rect 215 271 217 273
rect 256 271 258 273
rect 344 270 346 272
rect 394 270 396 272
rect 438 270 440 272
rect 494 270 496 272
rect 544 270 546 272
rect 594 270 596 272
rect 644 270 646 272
rect 103 238 105 240
rect 153 238 155 240
rect 224 239 226 241
rect 265 239 267 241
rect 353 238 355 240
rect 403 238 405 240
rect 447 238 449 240
rect 503 238 505 240
rect 553 238 555 240
rect 603 238 605 240
rect 653 238 655 240
rect 698 246 700 248
rect 717 246 719 248
rect 724 246 726 248
rect 798 246 800 248
rect 817 246 819 248
rect 824 246 826 248
rect 183 160 185 162
rect 104 152 106 154
rect 123 152 125 154
rect 130 152 132 154
rect 193 152 195 154
rect 233 152 235 154
rect 252 152 254 154
rect 259 152 261 154
rect 407 160 409 162
rect 328 152 330 154
rect 347 152 349 154
rect 354 152 356 154
rect 417 152 419 154
rect 457 152 459 154
rect 476 152 478 154
rect 483 152 485 154
rect 631 160 633 162
rect 552 152 554 154
rect 571 152 573 154
rect 578 152 580 154
rect 641 152 643 154
rect 766 176 768 178
rect 681 152 683 154
rect 700 152 702 154
rect 707 152 709 154
rect 775 144 777 146
rect 93 82 95 84
rect 226 66 228 68
rect 102 50 104 52
rect 147 58 149 60
rect 166 58 168 60
rect 173 58 175 60
rect 236 58 238 60
rect 360 82 362 84
rect 276 58 278 60
rect 295 58 297 60
rect 302 58 304 60
rect 492 66 494 68
rect 369 50 371 52
rect 413 58 415 60
rect 432 58 434 60
rect 439 58 441 60
rect 502 58 504 60
rect 627 82 629 84
rect 542 58 544 60
rect 561 58 563 60
rect 568 58 570 60
rect 758 66 760 68
rect 636 50 638 52
rect 679 58 681 60
rect 698 58 700 60
rect 705 58 707 60
rect 768 58 770 60
rect 892 82 894 84
rect 808 58 810 60
rect 827 58 829 60
rect 834 58 836 60
rect 901 50 903 52
<< ndifct0 >>
rect 87 320 89 322
rect 97 323 99 325
rect 107 331 109 333
rect 117 331 119 333
rect 117 324 119 326
rect 127 324 129 326
rect 144 317 146 319
rect 187 320 189 322
rect 197 323 199 325
rect 207 331 209 333
rect 217 331 219 333
rect 217 324 219 326
rect 227 324 229 326
rect 244 317 246 319
rect 276 326 278 328
rect 286 326 288 328
rect 296 326 298 328
rect 316 320 318 322
rect 326 323 328 325
rect 336 331 338 333
rect 346 331 348 333
rect 346 324 348 326
rect 356 324 358 326
rect 373 317 375 319
rect 411 320 413 322
rect 421 323 423 325
rect 431 331 433 333
rect 441 331 443 333
rect 441 324 443 326
rect 451 324 453 326
rect 468 317 470 319
rect 500 326 502 328
rect 510 326 512 328
rect 520 326 522 328
rect 540 320 542 322
rect 550 323 552 325
rect 560 331 562 333
rect 570 331 572 333
rect 570 324 572 326
rect 580 324 582 326
rect 597 317 599 319
rect 636 320 638 322
rect 646 323 648 325
rect 656 331 658 333
rect 666 331 668 333
rect 666 324 668 326
rect 676 324 678 326
rect 693 317 695 319
rect 754 323 756 325
rect 803 323 805 325
rect 853 323 855 325
rect 106 229 108 231
rect 156 229 158 231
rect 227 230 229 232
rect 268 230 270 232
rect 356 229 358 231
rect 406 229 408 231
rect 450 229 452 231
rect 506 229 508 231
rect 556 229 558 231
rect 606 229 608 231
rect 656 229 658 231
rect 681 226 683 228
rect 691 229 693 231
rect 701 237 703 239
rect 711 237 713 239
rect 711 230 713 232
rect 721 230 723 232
rect 738 223 740 225
rect 781 226 783 228
rect 791 229 793 231
rect 801 237 803 239
rect 811 237 813 239
rect 811 230 813 232
rect 821 230 823 232
rect 838 223 840 225
rect 87 132 89 134
rect 97 135 99 137
rect 107 143 109 145
rect 117 143 119 145
rect 117 136 119 138
rect 127 136 129 138
rect 144 129 146 131
rect 176 138 178 140
rect 186 138 188 140
rect 196 138 198 140
rect 216 132 218 134
rect 226 135 228 137
rect 236 143 238 145
rect 246 143 248 145
rect 246 136 248 138
rect 256 136 258 138
rect 273 129 275 131
rect 311 132 313 134
rect 321 135 323 137
rect 331 143 333 145
rect 341 143 343 145
rect 341 136 343 138
rect 351 136 353 138
rect 368 129 370 131
rect 400 138 402 140
rect 410 138 412 140
rect 420 138 422 140
rect 440 132 442 134
rect 450 135 452 137
rect 460 143 462 145
rect 470 143 472 145
rect 470 136 472 138
rect 480 136 482 138
rect 497 129 499 131
rect 535 132 537 134
rect 545 135 547 137
rect 555 143 557 145
rect 565 143 567 145
rect 565 136 567 138
rect 575 136 577 138
rect 592 129 594 131
rect 624 138 626 140
rect 634 138 636 140
rect 644 138 646 140
rect 664 132 666 134
rect 674 135 676 137
rect 684 143 686 145
rect 694 143 696 145
rect 694 136 696 138
rect 704 136 706 138
rect 721 129 723 131
rect 778 135 780 137
rect 105 41 107 43
rect 130 38 132 40
rect 140 41 142 43
rect 150 49 152 51
rect 160 49 162 51
rect 160 42 162 44
rect 170 42 172 44
rect 187 35 189 37
rect 219 44 221 46
rect 229 44 231 46
rect 239 44 241 46
rect 259 38 261 40
rect 269 41 271 43
rect 279 49 281 51
rect 289 49 291 51
rect 289 42 291 44
rect 299 42 301 44
rect 316 35 318 37
rect 372 41 374 43
rect 396 38 398 40
rect 406 41 408 43
rect 416 49 418 51
rect 426 49 428 51
rect 426 42 428 44
rect 436 42 438 44
rect 453 35 455 37
rect 485 44 487 46
rect 495 44 497 46
rect 505 44 507 46
rect 525 38 527 40
rect 535 41 537 43
rect 545 49 547 51
rect 555 49 557 51
rect 555 42 557 44
rect 565 42 567 44
rect 582 35 584 37
rect 639 41 641 43
rect 662 38 664 40
rect 672 41 674 43
rect 682 49 684 51
rect 692 49 694 51
rect 692 42 694 44
rect 702 42 704 44
rect 719 35 721 37
rect 751 44 753 46
rect 761 44 763 46
rect 771 44 773 46
rect 791 38 793 40
rect 801 41 803 43
rect 811 49 813 51
rect 821 49 823 51
rect 821 42 823 44
rect 831 42 833 44
rect 848 35 850 37
rect 904 41 906 43
<< ndifct1 >>
rect 77 324 79 326
rect 155 324 157 326
rect 177 324 179 326
rect 255 324 257 326
rect 266 326 268 328
rect 306 324 308 326
rect 384 324 386 326
rect 401 324 403 326
rect 479 324 481 326
rect 490 326 492 328
rect 530 324 532 326
rect 608 324 610 326
rect 626 324 628 326
rect 704 324 706 326
rect 725 326 727 328
rect 774 326 776 328
rect 824 326 826 328
rect 736 314 738 316
rect 785 314 787 316
rect 835 314 837 316
rect 77 232 79 234
rect 127 232 129 234
rect 198 233 200 235
rect 239 233 241 235
rect 327 232 329 234
rect 88 220 90 222
rect 138 220 140 222
rect 209 221 211 223
rect 250 221 252 223
rect 377 232 379 234
rect 421 232 423 234
rect 477 232 479 234
rect 527 232 529 234
rect 577 232 579 234
rect 627 232 629 234
rect 671 230 673 232
rect 338 220 340 222
rect 388 220 390 222
rect 432 220 434 222
rect 488 220 490 222
rect 538 220 540 222
rect 588 220 590 222
rect 638 220 640 222
rect 749 230 751 232
rect 771 230 773 232
rect 849 230 851 232
rect 77 136 79 138
rect 155 136 157 138
rect 166 138 168 140
rect 206 136 208 138
rect 284 136 286 138
rect 379 136 381 138
rect 390 138 392 140
rect 430 136 432 138
rect 508 136 510 138
rect 525 136 527 138
rect 603 136 605 138
rect 614 138 616 140
rect 654 136 656 138
rect 732 136 734 138
rect 749 138 751 140
rect 760 126 762 128
rect 76 44 78 46
rect 120 42 122 44
rect 87 32 89 34
rect 198 42 200 44
rect 209 44 211 46
rect 249 42 251 44
rect 327 42 329 44
rect 343 44 345 46
rect 386 42 388 44
rect 354 32 356 34
rect 464 42 466 44
rect 475 44 477 46
rect 515 42 517 44
rect 593 42 595 44
rect 610 44 612 46
rect 652 42 654 44
rect 621 32 623 34
rect 730 42 732 44
rect 741 44 743 46
rect 781 42 783 44
rect 859 42 861 44
rect 875 44 877 46
rect 886 32 888 34
<< ntiect1 >>
rect 267 374 269 376
rect 491 374 493 376
rect 726 374 728 376
rect 740 374 742 376
rect 754 374 756 376
rect 775 374 777 376
rect 789 374 791 376
rect 803 374 805 376
rect 825 374 827 376
rect 839 374 841 376
rect 853 374 855 376
rect 78 280 80 282
rect 92 280 94 282
rect 106 280 108 282
rect 128 280 130 282
rect 142 280 144 282
rect 156 280 158 282
rect 199 281 201 283
rect 213 281 215 283
rect 227 281 229 283
rect 240 281 242 283
rect 254 281 256 283
rect 268 281 270 283
rect 328 280 330 282
rect 342 280 344 282
rect 356 280 358 282
rect 378 280 380 282
rect 392 280 394 282
rect 406 280 408 282
rect 422 280 424 282
rect 436 280 438 282
rect 450 280 452 282
rect 478 280 480 282
rect 492 280 494 282
rect 506 280 508 282
rect 528 280 530 282
rect 542 280 544 282
rect 556 280 558 282
rect 578 280 580 282
rect 592 280 594 282
rect 606 280 608 282
rect 628 280 630 282
rect 642 280 644 282
rect 656 280 658 282
rect 167 186 169 188
rect 391 186 393 188
rect 615 186 617 188
rect 750 186 752 188
rect 764 186 766 188
rect 778 186 780 188
rect 77 92 79 94
rect 91 92 93 94
rect 105 92 107 94
rect 210 92 212 94
rect 344 92 346 94
rect 358 92 360 94
rect 372 92 374 94
rect 476 92 478 94
rect 611 92 613 94
rect 625 92 627 94
rect 639 92 641 94
rect 742 92 744 94
rect 876 92 878 94
rect 890 92 892 94
rect 904 92 906 94
<< ptiect1 >>
rect 267 314 269 316
rect 295 314 297 316
rect 491 314 493 316
rect 519 314 521 316
rect 726 314 728 316
rect 775 314 777 316
rect 825 314 827 316
rect 78 220 80 222
rect 128 220 130 222
rect 199 221 201 223
rect 240 221 242 223
rect 328 220 330 222
rect 378 220 380 222
rect 422 220 424 222
rect 478 220 480 222
rect 528 220 530 222
rect 578 220 580 222
rect 628 220 630 222
rect 167 126 169 128
rect 195 126 197 128
rect 391 126 393 128
rect 419 126 421 128
rect 615 126 617 128
rect 643 126 645 128
rect 750 126 752 128
rect 77 32 79 34
rect 238 32 240 34
rect 344 32 346 34
rect 504 32 506 34
rect 611 32 613 34
rect 770 32 772 34
rect 876 32 878 34
<< pdifct0 >>
rect 88 371 90 373
rect 100 352 102 354
rect 123 371 125 373
rect 123 364 125 366
rect 135 363 137 365
rect 135 356 137 358
rect 145 371 147 373
rect 145 364 147 366
rect 188 371 190 373
rect 200 352 202 354
rect 223 371 225 373
rect 223 364 225 366
rect 235 363 237 365
rect 235 356 237 358
rect 245 371 247 373
rect 245 364 247 366
rect 278 371 280 373
rect 296 364 298 366
rect 317 371 319 373
rect 329 352 331 354
rect 352 371 354 373
rect 352 364 354 366
rect 364 363 366 365
rect 364 356 366 358
rect 374 371 376 373
rect 374 364 376 366
rect 412 371 414 373
rect 424 352 426 354
rect 447 371 449 373
rect 447 364 449 366
rect 459 363 461 365
rect 459 356 461 358
rect 469 371 471 373
rect 469 364 471 366
rect 502 371 504 373
rect 520 364 522 366
rect 541 371 543 373
rect 553 352 555 354
rect 576 371 578 373
rect 576 364 578 366
rect 588 363 590 365
rect 588 356 590 358
rect 598 371 600 373
rect 598 364 600 366
rect 637 371 639 373
rect 649 352 651 354
rect 672 371 674 373
rect 672 364 674 366
rect 684 363 686 365
rect 684 356 686 358
rect 694 371 696 373
rect 694 364 696 366
rect 735 349 737 351
rect 745 349 747 351
rect 755 353 757 355
rect 784 349 786 351
rect 794 349 796 351
rect 804 353 806 355
rect 834 349 836 351
rect 844 349 846 351
rect 854 353 856 355
rect 87 255 89 257
rect 97 255 99 257
rect 107 259 109 261
rect 137 255 139 257
rect 147 255 149 257
rect 157 259 159 261
rect 208 256 210 258
rect 218 256 220 258
rect 228 260 230 262
rect 249 256 251 258
rect 259 256 261 258
rect 269 260 271 262
rect 337 255 339 257
rect 347 255 349 257
rect 357 259 359 261
rect 387 255 389 257
rect 397 255 399 257
rect 407 259 409 261
rect 431 255 433 257
rect 441 255 443 257
rect 451 259 453 261
rect 487 255 489 257
rect 497 255 499 257
rect 507 259 509 261
rect 537 255 539 257
rect 547 255 549 257
rect 557 259 559 261
rect 587 255 589 257
rect 597 255 599 257
rect 607 259 609 261
rect 637 255 639 257
rect 647 255 649 257
rect 657 259 659 261
rect 682 277 684 279
rect 694 258 696 260
rect 717 277 719 279
rect 717 270 719 272
rect 729 269 731 271
rect 729 262 731 264
rect 739 277 741 279
rect 739 270 741 272
rect 782 277 784 279
rect 794 258 796 260
rect 817 277 819 279
rect 817 270 819 272
rect 829 269 831 271
rect 829 262 831 264
rect 839 277 841 279
rect 839 270 841 272
rect 88 183 90 184
rect 100 164 102 166
rect 123 183 125 185
rect 123 176 125 178
rect 135 175 137 177
rect 135 168 137 170
rect 145 183 147 185
rect 145 176 147 178
rect 178 183 180 185
rect 196 176 198 178
rect 217 183 219 185
rect 229 164 231 166
rect 252 183 254 185
rect 252 176 254 178
rect 264 175 266 177
rect 264 168 266 170
rect 274 183 276 185
rect 274 176 276 178
rect 312 183 314 185
rect 324 164 326 166
rect 347 183 349 185
rect 347 176 349 178
rect 359 175 361 177
rect 359 168 361 170
rect 369 183 371 185
rect 369 176 371 178
rect 402 183 404 185
rect 420 176 422 178
rect 441 183 443 185
rect 453 164 455 166
rect 476 183 478 185
rect 476 176 478 178
rect 488 175 490 177
rect 488 168 490 170
rect 498 183 500 185
rect 498 176 500 178
rect 536 183 538 185
rect 548 164 550 166
rect 571 183 573 185
rect 571 176 573 178
rect 583 175 585 177
rect 583 168 585 170
rect 593 183 595 185
rect 593 176 595 178
rect 626 183 628 185
rect 644 176 646 178
rect 665 183 667 185
rect 677 164 679 166
rect 700 183 702 185
rect 700 176 702 178
rect 712 175 714 177
rect 712 168 714 170
rect 722 183 724 185
rect 722 176 724 178
rect 759 161 761 163
rect 769 161 771 163
rect 779 165 781 167
rect 86 67 88 69
rect 96 67 98 69
rect 106 71 108 73
rect 131 89 133 91
rect 143 70 145 72
rect 166 89 168 91
rect 166 82 168 84
rect 178 81 180 83
rect 178 74 180 76
rect 188 89 190 91
rect 188 82 190 84
rect 221 89 223 91
rect 239 82 241 84
rect 260 89 262 91
rect 272 70 274 72
rect 295 89 297 91
rect 295 82 297 84
rect 307 81 309 83
rect 307 74 309 76
rect 317 89 319 91
rect 317 82 319 84
rect 353 67 355 69
rect 363 67 365 69
rect 373 71 375 73
rect 397 89 399 91
rect 409 70 411 72
rect 432 89 434 91
rect 432 82 434 84
rect 444 81 446 83
rect 444 74 446 76
rect 454 89 456 91
rect 454 82 456 84
rect 487 89 489 91
rect 505 82 507 84
rect 526 89 528 91
rect 538 70 540 72
rect 561 89 563 91
rect 561 82 563 84
rect 573 81 575 83
rect 573 74 575 76
rect 583 89 585 91
rect 583 82 585 84
rect 620 67 622 69
rect 630 67 632 69
rect 640 71 642 73
rect 663 89 665 91
rect 675 70 677 72
rect 698 89 700 91
rect 698 82 700 84
rect 710 81 712 83
rect 710 74 712 76
rect 720 89 722 91
rect 720 82 722 84
rect 753 89 755 91
rect 771 82 773 84
rect 792 89 794 91
rect 804 70 806 72
rect 827 89 829 91
rect 827 82 829 84
rect 839 81 841 83
rect 839 74 841 76
rect 849 89 851 91
rect 849 82 851 84
rect 885 67 887 69
rect 895 67 897 69
rect 905 71 907 73
<< pdifct1 >>
rect 77 359 79 361
rect 77 352 79 354
rect 155 356 157 358
rect 155 349 157 351
rect 177 359 179 361
rect 177 352 179 354
rect 266 362 268 364
rect 255 356 257 358
rect 306 359 308 361
rect 255 349 257 351
rect 306 352 308 354
rect 384 356 386 358
rect 384 349 386 351
rect 401 359 403 361
rect 401 352 403 354
rect 490 362 492 364
rect 479 356 481 358
rect 530 359 532 361
rect 479 349 481 351
rect 530 352 532 354
rect 608 356 610 358
rect 608 349 610 351
rect 626 359 628 361
rect 626 352 628 354
rect 704 356 706 358
rect 704 349 706 351
rect 725 349 727 351
rect 774 349 776 351
rect 824 349 826 351
rect 77 255 79 257
rect 127 255 129 257
rect 198 256 200 258
rect 239 256 241 258
rect 327 255 329 257
rect 377 255 379 257
rect 421 255 423 257
rect 477 255 479 257
rect 527 255 529 257
rect 577 255 579 257
rect 627 255 629 257
rect 671 265 673 267
rect 671 258 673 260
rect 749 262 751 264
rect 749 255 751 257
rect 771 265 773 267
rect 771 258 773 260
rect 849 262 851 264
rect 849 255 851 257
rect 77 171 79 173
rect 77 164 79 166
rect 88 184 90 185
rect 166 174 168 176
rect 155 168 157 170
rect 206 171 208 173
rect 155 161 157 163
rect 206 164 208 166
rect 284 168 286 170
rect 284 161 286 163
rect 301 171 303 173
rect 301 164 303 166
rect 390 174 392 176
rect 379 168 381 170
rect 430 171 432 173
rect 379 161 381 163
rect 430 164 432 166
rect 508 168 510 170
rect 508 161 510 163
rect 525 171 527 173
rect 525 164 527 166
rect 614 174 616 176
rect 603 168 605 170
rect 654 171 656 173
rect 603 161 605 163
rect 654 164 656 166
rect 732 168 734 170
rect 732 161 734 163
rect 749 161 751 163
rect 76 67 78 69
rect 120 77 122 79
rect 120 70 122 72
rect 209 80 211 82
rect 198 74 200 76
rect 249 77 251 79
rect 198 67 200 69
rect 249 70 251 72
rect 327 74 329 76
rect 327 67 329 69
rect 343 67 345 69
rect 386 77 388 79
rect 386 70 388 72
rect 475 80 477 82
rect 464 74 466 76
rect 515 77 517 79
rect 464 67 466 69
rect 515 70 517 72
rect 593 74 595 76
rect 593 67 595 69
rect 610 67 612 69
rect 652 77 654 79
rect 652 70 654 72
rect 741 80 743 82
rect 730 74 732 76
rect 781 77 783 79
rect 730 67 732 69
rect 781 70 783 72
rect 859 74 861 76
rect 859 67 861 69
rect 875 67 877 69
<< alu0 >>
rect 86 371 88 373
rect 90 371 92 373
rect 86 370 92 371
rect 121 371 123 373
rect 125 371 127 373
rect 121 366 127 371
rect 143 371 145 373
rect 147 371 149 373
rect 121 364 123 366
rect 125 364 127 366
rect 121 363 127 364
rect 134 365 138 367
rect 134 363 135 365
rect 137 363 138 365
rect 143 366 149 371
rect 186 371 188 373
rect 190 371 192 373
rect 186 370 192 371
rect 221 371 223 373
rect 225 371 227 373
rect 143 364 145 366
rect 147 364 149 366
rect 143 363 149 364
rect 221 366 227 371
rect 243 371 245 373
rect 247 371 249 373
rect 221 364 223 366
rect 225 364 227 366
rect 221 363 227 364
rect 234 365 238 367
rect 234 363 235 365
rect 237 363 238 365
rect 243 366 249 371
rect 276 371 278 373
rect 280 371 282 373
rect 276 370 282 371
rect 315 371 317 373
rect 319 371 321 373
rect 315 370 321 371
rect 350 371 352 373
rect 354 371 356 373
rect 243 364 245 366
rect 247 364 249 366
rect 243 363 249 364
rect 91 359 115 363
rect 134 359 138 363
rect 89 355 95 359
rect 111 358 151 359
rect 111 356 135 358
rect 137 356 151 358
rect 89 345 93 355
rect 99 354 103 356
rect 111 355 151 356
rect 99 352 100 354
rect 102 352 103 354
rect 99 351 103 352
rect 89 343 90 345
rect 92 343 93 345
rect 89 341 93 343
rect 96 347 103 351
rect 96 336 100 347
rect 139 342 143 347
rect 139 340 140 342
rect 142 340 143 342
rect 82 335 100 336
rect 82 333 84 335
rect 86 334 100 335
rect 86 333 111 334
rect 82 332 107 333
rect 96 331 107 332
rect 109 331 111 333
rect 96 330 111 331
rect 116 333 120 335
rect 116 331 117 333
rect 119 331 120 333
rect 116 326 120 331
rect 139 338 143 340
rect 147 344 151 355
rect 147 342 153 344
rect 147 340 150 342
rect 152 340 153 342
rect 147 338 153 340
rect 147 335 151 338
rect 131 331 151 335
rect 131 327 135 331
rect 191 359 215 363
rect 234 359 238 363
rect 280 366 300 367
rect 280 364 296 366
rect 298 364 300 366
rect 280 363 300 364
rect 350 366 356 371
rect 372 371 374 373
rect 376 371 378 373
rect 350 364 352 366
rect 354 364 356 366
rect 350 363 356 364
rect 363 365 367 367
rect 363 363 364 365
rect 366 363 367 365
rect 372 366 378 371
rect 410 371 412 373
rect 414 371 416 373
rect 410 370 416 371
rect 445 371 447 373
rect 449 371 451 373
rect 372 364 374 366
rect 376 364 378 366
rect 372 363 378 364
rect 445 366 451 371
rect 467 371 469 373
rect 471 371 473 373
rect 445 364 447 366
rect 449 364 451 366
rect 445 363 451 364
rect 458 365 462 367
rect 458 363 459 365
rect 461 363 462 365
rect 467 366 473 371
rect 500 371 502 373
rect 504 371 506 373
rect 500 370 506 371
rect 539 371 541 373
rect 543 371 545 373
rect 539 370 545 371
rect 574 371 576 373
rect 578 371 580 373
rect 467 364 469 366
rect 471 364 473 366
rect 467 363 473 364
rect 189 355 195 359
rect 211 358 251 359
rect 211 356 235 358
rect 237 356 251 358
rect 189 345 193 355
rect 199 354 203 356
rect 211 355 251 356
rect 199 352 200 354
rect 202 352 203 354
rect 199 351 203 352
rect 189 343 190 345
rect 192 343 193 345
rect 189 341 193 343
rect 196 347 203 351
rect 196 336 200 347
rect 239 342 243 347
rect 239 340 240 342
rect 242 340 243 342
rect 182 335 200 336
rect 182 333 184 335
rect 186 334 200 335
rect 186 333 211 334
rect 182 332 207 333
rect 196 331 207 332
rect 209 331 211 333
rect 196 330 211 331
rect 216 333 220 335
rect 216 331 217 333
rect 219 331 220 333
rect 95 325 117 326
rect 86 322 90 324
rect 95 323 97 325
rect 99 324 117 325
rect 119 324 120 326
rect 99 323 120 324
rect 125 326 135 327
rect 125 324 127 326
rect 129 324 135 326
rect 125 323 135 324
rect 95 322 120 323
rect 216 326 220 331
rect 239 338 243 340
rect 247 344 251 355
rect 247 342 253 344
rect 247 340 250 342
rect 252 340 253 342
rect 247 338 253 340
rect 247 335 251 338
rect 231 331 251 335
rect 231 327 235 331
rect 195 325 217 326
rect 186 322 190 324
rect 195 323 197 325
rect 199 324 217 325
rect 219 324 220 326
rect 199 323 220 324
rect 225 326 235 327
rect 225 324 227 326
rect 229 324 235 326
rect 225 323 235 324
rect 268 360 269 363
rect 280 359 284 363
rect 272 355 284 359
rect 272 343 276 355
rect 320 359 344 363
rect 363 359 367 363
rect 272 341 273 343
rect 275 341 276 343
rect 272 336 276 341
rect 318 355 324 359
rect 340 358 380 359
rect 340 356 364 358
rect 366 356 380 358
rect 318 345 322 355
rect 328 354 332 356
rect 340 355 380 356
rect 328 352 329 354
rect 331 352 332 354
rect 328 351 332 352
rect 318 343 319 345
rect 321 343 322 345
rect 318 341 322 343
rect 325 347 332 351
rect 272 332 289 336
rect 195 322 220 323
rect 274 328 280 329
rect 274 326 276 328
rect 278 326 280 328
rect 86 320 87 322
rect 89 320 90 322
rect 186 320 187 322
rect 189 320 190 322
rect 86 317 90 320
rect 142 319 148 320
rect 142 317 144 319
rect 146 317 148 319
rect 186 317 190 320
rect 242 319 248 320
rect 242 317 244 319
rect 246 317 248 319
rect 274 317 280 326
rect 285 328 289 332
rect 285 326 286 328
rect 288 326 289 328
rect 285 324 289 326
rect 294 328 300 329
rect 294 326 296 328
rect 298 326 300 328
rect 294 317 300 326
rect 325 336 329 347
rect 368 342 372 347
rect 368 340 369 342
rect 371 340 372 342
rect 311 335 329 336
rect 311 333 313 335
rect 315 334 329 335
rect 315 333 340 334
rect 311 332 336 333
rect 325 331 336 332
rect 338 331 340 333
rect 325 330 340 331
rect 345 333 349 335
rect 345 331 346 333
rect 348 331 349 333
rect 345 326 349 331
rect 368 338 372 340
rect 376 344 380 355
rect 376 342 382 344
rect 376 340 379 342
rect 381 340 382 342
rect 376 338 382 340
rect 376 335 380 338
rect 360 331 380 335
rect 360 327 364 331
rect 324 325 346 326
rect 315 322 319 324
rect 324 323 326 325
rect 328 324 346 325
rect 348 324 349 326
rect 328 323 349 324
rect 354 326 364 327
rect 354 324 356 326
rect 358 324 364 326
rect 354 323 364 324
rect 415 359 439 363
rect 458 359 462 363
rect 504 366 524 367
rect 504 364 520 366
rect 522 364 524 366
rect 504 363 524 364
rect 574 366 580 371
rect 596 371 598 373
rect 600 371 602 373
rect 574 364 576 366
rect 578 364 580 366
rect 574 363 580 364
rect 587 365 591 367
rect 587 363 588 365
rect 590 363 591 365
rect 596 366 602 371
rect 635 371 637 373
rect 639 371 641 373
rect 635 370 641 371
rect 670 371 672 373
rect 674 371 676 373
rect 596 364 598 366
rect 600 364 602 366
rect 596 363 602 364
rect 670 366 676 371
rect 692 371 694 373
rect 696 371 698 373
rect 670 364 672 366
rect 674 364 676 366
rect 670 363 676 364
rect 683 365 687 367
rect 683 363 684 365
rect 686 363 687 365
rect 692 366 698 371
rect 692 364 694 366
rect 696 364 698 366
rect 692 363 698 364
rect 413 355 419 359
rect 435 358 475 359
rect 435 356 459 358
rect 461 356 475 358
rect 413 345 417 355
rect 423 354 427 356
rect 435 355 475 356
rect 423 352 424 354
rect 426 352 427 354
rect 423 351 427 352
rect 413 343 414 345
rect 416 343 417 345
rect 413 341 417 343
rect 420 347 427 351
rect 420 336 424 347
rect 463 342 467 347
rect 463 340 464 342
rect 466 340 467 342
rect 406 335 424 336
rect 406 333 408 335
rect 410 334 424 335
rect 410 333 435 334
rect 406 332 431 333
rect 420 331 431 332
rect 433 331 435 333
rect 420 330 435 331
rect 440 333 444 335
rect 440 331 441 333
rect 443 331 444 333
rect 440 326 444 331
rect 463 338 467 340
rect 471 344 475 355
rect 471 342 477 344
rect 471 340 474 342
rect 476 340 477 342
rect 471 338 477 340
rect 471 335 475 338
rect 455 331 475 335
rect 455 327 459 331
rect 419 325 441 326
rect 324 322 349 323
rect 410 322 414 324
rect 419 323 421 325
rect 423 324 441 325
rect 443 324 444 326
rect 423 323 444 324
rect 449 326 459 327
rect 449 324 451 326
rect 453 324 459 326
rect 449 323 459 324
rect 492 360 493 363
rect 504 359 508 363
rect 496 355 508 359
rect 496 343 500 355
rect 544 359 568 363
rect 587 359 591 363
rect 496 341 497 343
rect 499 341 500 343
rect 496 336 500 341
rect 542 355 548 359
rect 564 358 604 359
rect 564 356 588 358
rect 590 356 604 358
rect 542 345 546 355
rect 552 354 556 356
rect 564 355 604 356
rect 552 352 553 354
rect 555 352 556 354
rect 552 351 556 352
rect 542 343 543 345
rect 545 343 546 345
rect 542 341 546 343
rect 549 347 556 351
rect 496 332 513 336
rect 419 322 444 323
rect 498 328 504 329
rect 498 326 500 328
rect 502 326 504 328
rect 315 320 316 322
rect 318 320 319 322
rect 410 320 411 322
rect 413 320 414 322
rect 315 317 319 320
rect 371 319 377 320
rect 371 317 373 319
rect 375 317 377 319
rect 410 317 414 320
rect 466 319 472 320
rect 466 317 468 319
rect 470 317 472 319
rect 498 317 504 326
rect 509 328 513 332
rect 509 326 510 328
rect 512 326 513 328
rect 509 324 513 326
rect 518 328 524 329
rect 518 326 520 328
rect 522 326 524 328
rect 518 317 524 326
rect 549 336 553 347
rect 592 342 596 347
rect 592 340 593 342
rect 595 340 596 342
rect 535 335 553 336
rect 535 333 537 335
rect 539 334 553 335
rect 539 333 564 334
rect 535 332 560 333
rect 549 331 560 332
rect 562 331 564 333
rect 549 330 564 331
rect 569 333 573 335
rect 569 331 570 333
rect 572 331 573 333
rect 569 326 573 331
rect 592 338 596 340
rect 600 344 604 355
rect 600 342 606 344
rect 600 340 603 342
rect 605 340 606 342
rect 600 338 606 340
rect 600 335 604 338
rect 584 331 604 335
rect 584 327 588 331
rect 548 325 570 326
rect 539 322 543 324
rect 548 323 550 325
rect 552 324 570 325
rect 572 324 573 326
rect 552 323 573 324
rect 578 326 588 327
rect 578 324 580 326
rect 582 324 588 326
rect 578 323 588 324
rect 640 359 664 363
rect 683 359 687 363
rect 638 355 644 359
rect 660 358 700 359
rect 660 356 684 358
rect 686 356 700 358
rect 638 345 642 355
rect 648 354 652 356
rect 660 355 700 356
rect 648 352 649 354
rect 651 352 652 354
rect 648 351 652 352
rect 638 343 639 345
rect 641 343 642 345
rect 638 341 642 343
rect 645 347 652 351
rect 645 336 649 347
rect 688 342 692 347
rect 688 340 689 342
rect 691 340 692 342
rect 631 335 649 336
rect 688 338 692 340
rect 696 344 700 355
rect 696 342 702 344
rect 696 340 699 342
rect 701 340 702 342
rect 696 338 702 340
rect 696 335 700 338
rect 631 333 633 335
rect 635 334 649 335
rect 635 333 660 334
rect 631 332 656 333
rect 645 331 656 332
rect 658 331 660 333
rect 645 330 660 331
rect 665 333 669 335
rect 665 331 666 333
rect 668 331 669 333
rect 665 326 669 331
rect 680 331 700 335
rect 680 327 684 331
rect 644 325 666 326
rect 548 322 573 323
rect 635 322 639 324
rect 644 323 646 325
rect 648 324 666 325
rect 668 324 669 326
rect 648 323 669 324
rect 674 326 684 327
rect 674 324 676 326
rect 678 324 684 326
rect 674 323 684 324
rect 727 347 728 353
rect 731 352 735 373
rect 754 355 758 373
rect 754 353 755 355
rect 757 353 758 355
rect 731 351 739 352
rect 731 349 735 351
rect 737 349 739 351
rect 731 348 739 349
rect 743 351 749 352
rect 754 351 758 353
rect 743 349 745 351
rect 747 349 749 351
rect 743 343 749 349
rect 730 342 749 343
rect 730 340 732 342
rect 734 340 749 342
rect 730 339 749 340
rect 727 328 728 330
rect 644 322 669 323
rect 739 326 743 339
rect 776 347 777 353
rect 780 352 784 373
rect 803 355 807 373
rect 803 353 804 355
rect 806 353 807 355
rect 780 351 788 352
rect 780 349 784 351
rect 786 349 788 351
rect 780 348 788 349
rect 792 351 798 352
rect 803 351 807 353
rect 792 349 794 351
rect 796 349 798 351
rect 792 343 798 349
rect 779 342 798 343
rect 779 340 781 342
rect 783 340 798 342
rect 779 339 798 340
rect 776 328 777 330
rect 739 325 758 326
rect 739 323 754 325
rect 756 323 758 325
rect 739 322 758 323
rect 788 326 792 339
rect 826 347 827 353
rect 830 352 834 373
rect 853 355 857 373
rect 853 353 854 355
rect 856 353 857 355
rect 830 351 838 352
rect 830 349 834 351
rect 836 349 838 351
rect 830 348 838 349
rect 842 351 848 352
rect 853 351 857 353
rect 842 349 844 351
rect 846 349 848 351
rect 842 343 848 349
rect 829 342 848 343
rect 829 340 831 342
rect 833 340 848 342
rect 829 339 848 340
rect 826 328 827 330
rect 788 325 807 326
rect 788 323 803 325
rect 805 323 807 325
rect 788 322 807 323
rect 838 326 842 339
rect 838 325 857 326
rect 838 323 853 325
rect 855 323 857 325
rect 838 322 857 323
rect 539 320 540 322
rect 542 320 543 322
rect 635 320 636 322
rect 638 320 639 322
rect 539 317 543 320
rect 595 319 601 320
rect 595 317 597 319
rect 599 317 601 319
rect 635 317 639 320
rect 691 319 697 320
rect 691 317 693 319
rect 695 317 697 319
rect 79 253 80 259
rect 83 258 87 279
rect 106 261 110 279
rect 106 259 107 261
rect 109 259 110 261
rect 83 257 91 258
rect 83 255 87 257
rect 89 255 91 257
rect 83 254 91 255
rect 95 257 101 258
rect 106 257 110 259
rect 95 255 97 257
rect 99 255 101 257
rect 95 249 101 255
rect 82 248 101 249
rect 82 246 84 248
rect 86 246 101 248
rect 82 245 101 246
rect 79 234 80 236
rect 91 232 95 245
rect 129 253 130 259
rect 133 258 137 279
rect 156 261 160 279
rect 156 259 157 261
rect 159 259 160 261
rect 133 257 141 258
rect 133 255 137 257
rect 139 255 141 257
rect 133 254 141 255
rect 145 257 151 258
rect 156 257 160 259
rect 145 255 147 257
rect 149 255 151 257
rect 145 249 151 255
rect 132 248 151 249
rect 132 246 134 248
rect 136 246 151 248
rect 132 245 151 246
rect 129 234 130 236
rect 91 231 110 232
rect 91 229 106 231
rect 108 229 110 231
rect 91 228 110 229
rect 141 232 145 245
rect 200 254 201 260
rect 204 259 208 280
rect 227 262 231 280
rect 227 260 228 262
rect 230 260 231 262
rect 204 258 212 259
rect 204 256 208 258
rect 210 256 212 258
rect 204 255 212 256
rect 216 258 222 259
rect 227 258 231 260
rect 216 256 218 258
rect 220 256 222 258
rect 216 250 222 256
rect 203 249 222 250
rect 203 247 205 249
rect 207 247 222 249
rect 203 246 222 247
rect 200 235 201 237
rect 141 231 160 232
rect 141 229 156 231
rect 158 229 160 231
rect 212 233 216 246
rect 241 254 242 260
rect 245 259 249 280
rect 268 262 272 280
rect 268 260 269 262
rect 271 260 272 262
rect 245 258 253 259
rect 245 256 249 258
rect 251 256 253 258
rect 245 255 253 256
rect 257 258 263 259
rect 268 258 272 260
rect 257 256 259 258
rect 261 256 263 258
rect 257 250 263 256
rect 244 249 263 250
rect 244 247 246 249
rect 248 247 263 249
rect 244 246 263 247
rect 241 235 242 237
rect 212 232 231 233
rect 212 230 227 232
rect 229 230 231 232
rect 212 229 231 230
rect 253 233 257 246
rect 329 253 330 259
rect 333 258 337 279
rect 356 261 360 279
rect 356 259 357 261
rect 359 259 360 261
rect 333 257 341 258
rect 333 255 337 257
rect 339 255 341 257
rect 333 254 341 255
rect 345 257 351 258
rect 356 257 360 259
rect 345 255 347 257
rect 349 255 351 257
rect 345 249 351 255
rect 332 248 351 249
rect 332 246 334 248
rect 336 246 351 248
rect 332 245 351 246
rect 329 234 330 236
rect 253 232 272 233
rect 253 230 268 232
rect 270 230 272 232
rect 253 229 272 230
rect 141 228 160 229
rect 341 232 345 245
rect 379 253 380 259
rect 383 258 387 279
rect 406 261 410 279
rect 406 259 407 261
rect 409 259 410 261
rect 383 257 391 258
rect 383 255 387 257
rect 389 255 391 257
rect 383 254 391 255
rect 395 257 401 258
rect 406 257 410 259
rect 395 255 397 257
rect 399 255 401 257
rect 395 249 401 255
rect 382 248 401 249
rect 382 246 384 248
rect 386 246 401 248
rect 382 245 401 246
rect 379 234 380 236
rect 341 231 360 232
rect 341 229 356 231
rect 358 229 360 231
rect 341 228 360 229
rect 391 232 395 245
rect 423 253 424 259
rect 427 258 431 279
rect 450 261 454 279
rect 450 259 451 261
rect 453 259 454 261
rect 427 257 435 258
rect 427 255 431 257
rect 433 255 435 257
rect 427 254 435 255
rect 439 257 445 258
rect 450 257 454 259
rect 439 255 441 257
rect 443 255 445 257
rect 439 249 445 255
rect 426 248 445 249
rect 426 246 428 248
rect 430 246 445 248
rect 426 245 445 246
rect 423 234 424 236
rect 391 231 410 232
rect 391 229 406 231
rect 408 229 410 231
rect 391 228 410 229
rect 435 232 439 245
rect 479 253 480 259
rect 483 258 487 279
rect 506 261 510 279
rect 506 259 507 261
rect 509 259 510 261
rect 483 257 491 258
rect 483 255 487 257
rect 489 255 491 257
rect 483 254 491 255
rect 495 257 501 258
rect 506 257 510 259
rect 495 255 497 257
rect 499 255 501 257
rect 495 249 501 255
rect 482 248 501 249
rect 482 246 484 248
rect 486 246 501 248
rect 482 245 501 246
rect 479 234 480 236
rect 435 231 454 232
rect 435 229 450 231
rect 452 229 454 231
rect 435 228 454 229
rect 491 232 495 245
rect 529 253 530 259
rect 533 258 537 279
rect 556 261 560 279
rect 556 259 557 261
rect 559 259 560 261
rect 533 257 541 258
rect 533 255 537 257
rect 539 255 541 257
rect 533 254 541 255
rect 545 257 551 258
rect 556 257 560 259
rect 545 255 547 257
rect 549 255 551 257
rect 545 249 551 255
rect 532 248 551 249
rect 532 246 534 248
rect 536 246 551 248
rect 532 245 551 246
rect 529 234 530 236
rect 491 231 510 232
rect 491 229 506 231
rect 508 229 510 231
rect 491 228 510 229
rect 541 232 545 245
rect 579 253 580 259
rect 583 258 587 279
rect 606 261 610 279
rect 606 259 607 261
rect 609 259 610 261
rect 583 257 591 258
rect 583 255 587 257
rect 589 255 591 257
rect 583 254 591 255
rect 595 257 601 258
rect 606 257 610 259
rect 595 255 597 257
rect 599 255 601 257
rect 595 249 601 255
rect 582 248 601 249
rect 582 246 584 248
rect 586 246 601 248
rect 582 245 601 246
rect 579 234 580 236
rect 541 231 560 232
rect 541 229 556 231
rect 558 229 560 231
rect 541 228 560 229
rect 591 232 595 245
rect 629 253 630 259
rect 633 258 637 279
rect 656 261 660 279
rect 680 277 682 279
rect 684 277 686 279
rect 680 276 686 277
rect 715 277 717 279
rect 719 277 721 279
rect 656 259 657 261
rect 659 259 660 261
rect 633 257 641 258
rect 633 255 637 257
rect 639 255 641 257
rect 633 254 641 255
rect 645 257 651 258
rect 656 257 660 259
rect 715 272 721 277
rect 737 277 739 279
rect 741 277 743 279
rect 715 270 717 272
rect 719 270 721 272
rect 715 269 721 270
rect 728 271 732 273
rect 728 269 729 271
rect 731 269 732 271
rect 737 272 743 277
rect 780 277 782 279
rect 784 277 786 279
rect 780 276 786 277
rect 815 277 817 279
rect 819 277 821 279
rect 737 270 739 272
rect 741 270 743 272
rect 737 269 743 270
rect 815 272 821 277
rect 837 277 839 279
rect 841 277 843 279
rect 815 270 817 272
rect 819 270 821 272
rect 815 269 821 270
rect 828 271 832 273
rect 828 269 829 271
rect 831 269 832 271
rect 837 272 843 277
rect 837 270 839 272
rect 841 270 843 272
rect 837 269 843 270
rect 685 265 709 269
rect 728 265 732 269
rect 645 255 647 257
rect 649 255 651 257
rect 645 249 651 255
rect 683 261 689 265
rect 705 264 745 265
rect 705 262 729 264
rect 731 262 745 264
rect 632 248 651 249
rect 632 246 634 248
rect 636 246 651 248
rect 632 245 651 246
rect 629 234 630 236
rect 591 231 610 232
rect 591 229 606 231
rect 608 229 610 231
rect 591 228 610 229
rect 641 232 645 245
rect 683 251 687 261
rect 693 260 697 262
rect 705 261 745 262
rect 693 258 694 260
rect 696 258 697 260
rect 693 257 697 258
rect 683 249 684 251
rect 686 249 687 251
rect 683 247 687 249
rect 690 253 697 257
rect 690 242 694 253
rect 733 248 737 253
rect 733 246 734 248
rect 736 246 737 248
rect 676 241 694 242
rect 676 239 678 241
rect 680 240 694 241
rect 680 239 705 240
rect 676 238 701 239
rect 690 237 701 238
rect 703 237 705 239
rect 690 236 705 237
rect 710 239 714 241
rect 710 237 711 239
rect 713 237 714 239
rect 710 232 714 237
rect 733 244 737 246
rect 741 250 745 261
rect 741 248 747 250
rect 741 246 744 248
rect 746 246 747 248
rect 741 244 747 246
rect 741 241 745 244
rect 725 237 745 241
rect 725 233 729 237
rect 641 231 660 232
rect 641 229 656 231
rect 658 229 660 231
rect 641 228 660 229
rect 689 231 711 232
rect 680 228 684 230
rect 689 229 691 231
rect 693 230 711 231
rect 713 230 714 232
rect 693 229 714 230
rect 719 232 729 233
rect 719 230 721 232
rect 723 230 729 232
rect 719 229 729 230
rect 785 265 809 269
rect 828 265 832 269
rect 783 261 789 265
rect 805 264 845 265
rect 805 262 829 264
rect 831 262 845 264
rect 783 251 787 261
rect 793 260 797 262
rect 805 261 845 262
rect 793 258 794 260
rect 796 258 797 260
rect 793 257 797 258
rect 783 249 784 251
rect 786 249 787 251
rect 783 247 787 249
rect 790 253 797 257
rect 790 242 794 253
rect 833 248 837 253
rect 833 246 834 248
rect 836 246 837 248
rect 776 241 794 242
rect 776 239 778 241
rect 780 240 794 241
rect 780 239 805 240
rect 776 238 801 239
rect 790 237 801 238
rect 803 237 805 239
rect 790 236 805 237
rect 810 239 814 241
rect 810 237 811 239
rect 813 237 814 239
rect 810 232 814 237
rect 833 244 837 246
rect 841 250 845 261
rect 841 248 847 250
rect 841 246 844 248
rect 846 246 847 248
rect 841 244 847 246
rect 841 241 845 244
rect 825 237 845 241
rect 825 233 829 237
rect 789 231 811 232
rect 689 228 714 229
rect 780 228 784 230
rect 789 229 791 231
rect 793 230 811 231
rect 813 230 814 232
rect 793 229 814 230
rect 819 232 829 233
rect 819 230 821 232
rect 823 230 829 232
rect 819 229 829 230
rect 789 228 814 229
rect 680 226 681 228
rect 683 226 684 228
rect 780 226 781 228
rect 783 226 784 228
rect 680 223 684 226
rect 736 225 742 226
rect 736 223 738 225
rect 740 223 742 225
rect 780 223 784 226
rect 836 225 842 226
rect 836 223 838 225
rect 840 223 842 225
rect 86 183 88 184
rect 90 183 92 184
rect 86 182 92 183
rect 121 183 123 185
rect 125 183 127 185
rect 121 178 127 183
rect 143 183 145 185
rect 147 183 149 185
rect 121 176 123 178
rect 125 176 127 178
rect 121 175 127 176
rect 134 177 138 179
rect 134 175 135 177
rect 137 175 138 177
rect 143 178 149 183
rect 176 183 178 185
rect 180 183 182 185
rect 176 182 182 183
rect 215 183 217 185
rect 219 183 221 185
rect 215 182 221 183
rect 250 183 252 185
rect 254 183 256 185
rect 143 176 145 178
rect 147 176 149 178
rect 143 175 149 176
rect 91 171 115 175
rect 134 171 138 175
rect 180 178 200 179
rect 180 176 196 178
rect 198 176 200 178
rect 180 175 200 176
rect 250 178 256 183
rect 272 183 274 185
rect 276 183 278 185
rect 250 176 252 178
rect 254 176 256 178
rect 250 175 256 176
rect 263 177 267 179
rect 263 175 264 177
rect 266 175 267 177
rect 272 178 278 183
rect 310 183 312 185
rect 314 183 316 185
rect 310 182 316 183
rect 345 183 347 185
rect 349 183 351 185
rect 272 176 274 178
rect 276 176 278 178
rect 272 175 278 176
rect 345 178 351 183
rect 367 183 369 185
rect 371 183 373 185
rect 345 176 347 178
rect 349 176 351 178
rect 345 175 351 176
rect 358 177 362 179
rect 358 175 359 177
rect 361 175 362 177
rect 367 178 373 183
rect 400 183 402 185
rect 404 183 406 185
rect 400 182 406 183
rect 439 183 441 185
rect 443 183 445 185
rect 439 182 445 183
rect 474 183 476 185
rect 478 183 480 185
rect 367 176 369 178
rect 371 176 373 178
rect 367 175 373 176
rect 89 167 95 171
rect 111 170 151 171
rect 111 168 135 170
rect 137 168 151 170
rect 89 157 93 167
rect 99 166 103 168
rect 111 167 151 168
rect 99 164 100 166
rect 102 164 103 166
rect 99 163 103 164
rect 89 155 90 157
rect 92 155 93 157
rect 89 153 93 155
rect 96 159 103 163
rect 96 148 100 159
rect 139 154 143 159
rect 139 152 140 154
rect 142 152 143 154
rect 82 147 100 148
rect 82 145 84 147
rect 86 146 100 147
rect 86 145 111 146
rect 82 144 107 145
rect 96 143 107 144
rect 109 143 111 145
rect 96 142 111 143
rect 116 145 120 147
rect 116 143 117 145
rect 119 143 120 145
rect 116 138 120 143
rect 139 150 143 152
rect 147 156 151 167
rect 147 154 153 156
rect 147 152 150 154
rect 152 152 153 154
rect 147 150 153 152
rect 147 147 151 150
rect 131 143 151 147
rect 131 139 135 143
rect 95 137 117 138
rect 86 134 90 136
rect 95 135 97 137
rect 99 136 117 137
rect 119 136 120 138
rect 99 135 120 136
rect 125 138 135 139
rect 125 136 127 138
rect 129 136 135 138
rect 125 135 135 136
rect 168 172 169 175
rect 180 171 184 175
rect 172 167 184 171
rect 172 155 176 167
rect 220 171 244 175
rect 263 171 267 175
rect 172 153 173 155
rect 175 153 176 155
rect 172 148 176 153
rect 218 167 224 171
rect 240 170 280 171
rect 240 168 264 170
rect 266 168 280 170
rect 218 157 222 167
rect 228 166 232 168
rect 240 167 280 168
rect 228 164 229 166
rect 231 164 232 166
rect 228 163 232 164
rect 218 155 219 157
rect 221 155 222 157
rect 218 153 222 155
rect 225 159 232 163
rect 172 144 189 148
rect 95 134 120 135
rect 174 140 180 141
rect 174 138 176 140
rect 178 138 180 140
rect 86 132 87 134
rect 89 132 90 134
rect 86 129 90 132
rect 142 131 148 132
rect 142 129 144 131
rect 146 129 148 131
rect 174 129 180 138
rect 185 140 189 144
rect 185 138 186 140
rect 188 138 189 140
rect 185 136 189 138
rect 194 140 200 141
rect 194 138 196 140
rect 198 138 200 140
rect 194 129 200 138
rect 225 148 229 159
rect 268 154 272 159
rect 268 152 269 154
rect 271 152 272 154
rect 211 147 229 148
rect 268 150 272 152
rect 276 156 280 167
rect 276 154 282 156
rect 276 152 279 154
rect 281 152 282 154
rect 276 150 282 152
rect 211 145 213 147
rect 215 146 229 147
rect 215 145 240 146
rect 211 144 236 145
rect 225 143 236 144
rect 238 143 240 145
rect 225 142 240 143
rect 245 145 249 147
rect 245 143 246 145
rect 248 143 249 145
rect 245 138 249 143
rect 276 147 280 150
rect 260 143 280 147
rect 260 139 264 143
rect 315 171 339 175
rect 358 171 362 175
rect 404 178 424 179
rect 404 176 420 178
rect 422 176 424 178
rect 404 175 424 176
rect 474 178 480 183
rect 496 183 498 185
rect 500 183 502 185
rect 474 176 476 178
rect 478 176 480 178
rect 474 175 480 176
rect 487 177 491 179
rect 487 175 488 177
rect 490 175 491 177
rect 496 178 502 183
rect 534 183 536 185
rect 538 183 540 185
rect 534 182 540 183
rect 569 183 571 185
rect 573 183 575 185
rect 496 176 498 178
rect 500 176 502 178
rect 496 175 502 176
rect 569 178 575 183
rect 591 183 593 185
rect 595 183 597 185
rect 569 176 571 178
rect 573 176 575 178
rect 569 175 575 176
rect 582 177 586 179
rect 582 175 583 177
rect 585 175 586 177
rect 591 178 597 183
rect 624 183 626 185
rect 628 183 630 185
rect 624 182 630 183
rect 663 183 665 185
rect 667 183 669 185
rect 663 182 669 183
rect 698 183 700 185
rect 702 183 704 185
rect 591 176 593 178
rect 595 176 597 178
rect 591 175 597 176
rect 313 167 319 171
rect 335 170 375 171
rect 335 168 359 170
rect 361 168 375 170
rect 313 157 317 167
rect 323 166 327 168
rect 335 167 375 168
rect 323 164 324 166
rect 326 164 327 166
rect 323 163 327 164
rect 313 155 314 157
rect 316 155 317 157
rect 313 153 317 155
rect 320 159 327 163
rect 320 148 324 159
rect 363 154 367 159
rect 363 152 364 154
rect 366 152 367 154
rect 224 137 246 138
rect 215 134 219 136
rect 224 135 226 137
rect 228 136 246 137
rect 248 136 249 138
rect 228 135 249 136
rect 254 138 264 139
rect 254 136 256 138
rect 258 136 264 138
rect 254 135 264 136
rect 306 147 324 148
rect 306 145 308 147
rect 310 146 324 147
rect 310 145 335 146
rect 306 144 331 145
rect 320 143 331 144
rect 333 143 335 145
rect 320 142 335 143
rect 340 145 344 147
rect 340 143 341 145
rect 343 143 344 145
rect 224 134 249 135
rect 340 138 344 143
rect 363 150 367 152
rect 371 156 375 167
rect 371 154 377 156
rect 371 152 374 154
rect 376 152 377 154
rect 371 150 377 152
rect 371 147 375 150
rect 355 143 375 147
rect 355 139 359 143
rect 319 137 341 138
rect 310 134 314 136
rect 319 135 321 137
rect 323 136 341 137
rect 343 136 344 138
rect 323 135 344 136
rect 349 138 359 139
rect 349 136 351 138
rect 353 136 359 138
rect 349 135 359 136
rect 392 172 393 175
rect 404 171 408 175
rect 396 167 408 171
rect 396 155 400 167
rect 444 171 468 175
rect 487 171 491 175
rect 396 153 397 155
rect 399 153 400 155
rect 396 148 400 153
rect 442 167 448 171
rect 464 170 504 171
rect 464 168 488 170
rect 490 168 504 170
rect 442 157 446 167
rect 452 166 456 168
rect 464 167 504 168
rect 452 164 453 166
rect 455 164 456 166
rect 452 163 456 164
rect 442 155 443 157
rect 445 155 446 157
rect 442 153 446 155
rect 449 159 456 163
rect 396 144 413 148
rect 319 134 344 135
rect 398 140 404 141
rect 398 138 400 140
rect 402 138 404 140
rect 215 132 216 134
rect 218 132 219 134
rect 310 132 311 134
rect 313 132 314 134
rect 215 129 219 132
rect 271 131 277 132
rect 271 129 273 131
rect 275 129 277 131
rect 310 129 314 132
rect 366 131 372 132
rect 366 129 368 131
rect 370 129 372 131
rect 398 129 404 138
rect 409 140 413 144
rect 409 138 410 140
rect 412 138 413 140
rect 409 136 413 138
rect 418 140 424 141
rect 418 138 420 140
rect 422 138 424 140
rect 418 129 424 138
rect 449 148 453 159
rect 492 154 496 159
rect 492 152 493 154
rect 495 152 496 154
rect 435 147 453 148
rect 492 150 496 152
rect 500 156 504 167
rect 500 154 506 156
rect 500 152 503 154
rect 505 152 506 154
rect 500 150 506 152
rect 435 145 437 147
rect 439 146 453 147
rect 439 145 464 146
rect 435 144 460 145
rect 449 143 460 144
rect 462 143 464 145
rect 449 142 464 143
rect 469 145 473 147
rect 469 143 470 145
rect 472 143 473 145
rect 469 138 473 143
rect 500 147 504 150
rect 484 143 504 147
rect 484 139 488 143
rect 448 137 470 138
rect 439 134 443 136
rect 448 135 450 137
rect 452 136 470 137
rect 472 136 473 138
rect 452 135 473 136
rect 478 138 488 139
rect 478 136 480 138
rect 482 136 488 138
rect 478 135 488 136
rect 539 171 563 175
rect 582 171 586 175
rect 628 178 648 179
rect 628 176 644 178
rect 646 176 648 178
rect 628 175 648 176
rect 698 178 704 183
rect 720 183 722 185
rect 724 183 726 185
rect 698 176 700 178
rect 702 176 704 178
rect 698 175 704 176
rect 711 177 715 179
rect 711 175 712 177
rect 714 175 715 177
rect 720 178 726 183
rect 720 176 722 178
rect 724 176 726 178
rect 720 175 726 176
rect 537 167 543 171
rect 559 170 599 171
rect 559 168 583 170
rect 585 168 599 170
rect 537 157 541 167
rect 547 166 551 168
rect 559 167 599 168
rect 547 164 548 166
rect 550 164 551 166
rect 547 163 551 164
rect 537 155 538 157
rect 540 155 541 157
rect 537 153 541 155
rect 544 159 551 163
rect 544 148 548 159
rect 587 154 591 159
rect 587 152 588 154
rect 590 152 591 154
rect 530 147 548 148
rect 530 145 532 147
rect 534 146 548 147
rect 534 145 559 146
rect 530 144 555 145
rect 544 143 555 144
rect 557 143 559 145
rect 544 142 559 143
rect 564 145 568 147
rect 564 143 565 145
rect 567 143 568 145
rect 564 138 568 143
rect 587 150 591 152
rect 595 156 599 167
rect 595 154 601 156
rect 595 152 598 154
rect 600 152 601 154
rect 595 150 601 152
rect 595 147 599 150
rect 579 143 599 147
rect 579 139 583 143
rect 543 137 565 138
rect 448 134 473 135
rect 534 134 538 136
rect 543 135 545 137
rect 547 136 565 137
rect 567 136 568 138
rect 547 135 568 136
rect 573 138 583 139
rect 573 136 575 138
rect 577 136 583 138
rect 573 135 583 136
rect 616 172 617 175
rect 628 171 632 175
rect 620 167 632 171
rect 620 155 624 167
rect 668 171 692 175
rect 711 171 715 175
rect 620 153 621 155
rect 623 153 624 155
rect 620 148 624 153
rect 666 167 672 171
rect 688 170 728 171
rect 688 168 712 170
rect 714 168 728 170
rect 666 157 670 167
rect 676 166 680 168
rect 688 167 728 168
rect 676 164 677 166
rect 679 164 680 166
rect 676 163 680 164
rect 666 155 667 157
rect 669 155 670 157
rect 666 153 670 155
rect 673 159 680 163
rect 620 144 637 148
rect 543 134 568 135
rect 622 140 628 141
rect 622 138 624 140
rect 626 138 628 140
rect 439 132 440 134
rect 442 132 443 134
rect 534 132 535 134
rect 537 132 538 134
rect 439 129 443 132
rect 495 131 501 132
rect 495 129 497 131
rect 499 129 501 131
rect 534 129 538 132
rect 590 131 596 132
rect 590 129 592 131
rect 594 129 596 131
rect 622 129 628 138
rect 633 140 637 144
rect 633 138 634 140
rect 636 138 637 140
rect 633 136 637 138
rect 642 140 648 141
rect 642 138 644 140
rect 646 138 648 140
rect 642 129 648 138
rect 673 148 677 159
rect 716 154 720 159
rect 716 152 717 154
rect 719 152 720 154
rect 659 147 677 148
rect 659 145 661 147
rect 663 146 677 147
rect 663 145 688 146
rect 659 144 684 145
rect 673 143 684 144
rect 686 143 688 145
rect 673 142 688 143
rect 693 145 697 147
rect 693 143 694 145
rect 696 143 697 145
rect 693 138 697 143
rect 716 150 720 152
rect 724 156 728 167
rect 724 154 730 156
rect 724 152 727 154
rect 729 152 730 154
rect 724 150 730 152
rect 724 147 728 150
rect 708 143 728 147
rect 708 139 712 143
rect 672 137 694 138
rect 663 134 667 136
rect 672 135 674 137
rect 676 136 694 137
rect 696 136 697 138
rect 676 135 697 136
rect 702 138 712 139
rect 702 136 704 138
rect 706 136 712 138
rect 702 135 712 136
rect 751 159 752 165
rect 755 164 759 185
rect 778 167 782 185
rect 778 165 779 167
rect 781 165 782 167
rect 755 163 763 164
rect 755 161 759 163
rect 761 161 763 163
rect 755 160 763 161
rect 767 163 773 164
rect 778 163 782 165
rect 767 161 769 163
rect 771 161 773 163
rect 767 155 773 161
rect 754 154 773 155
rect 754 152 756 154
rect 758 152 773 154
rect 754 151 773 152
rect 751 140 752 142
rect 672 134 697 135
rect 763 138 767 151
rect 763 137 782 138
rect 763 135 778 137
rect 780 135 782 137
rect 763 134 782 135
rect 663 132 664 134
rect 666 132 667 134
rect 663 129 667 132
rect 719 131 725 132
rect 719 129 721 131
rect 723 129 725 131
rect 78 65 79 71
rect 82 70 86 91
rect 105 73 109 91
rect 129 89 131 91
rect 133 89 135 91
rect 129 88 135 89
rect 164 89 166 91
rect 168 89 170 91
rect 105 71 106 73
rect 108 71 109 73
rect 82 69 90 70
rect 82 67 86 69
rect 88 67 90 69
rect 82 66 90 67
rect 94 69 100 70
rect 105 69 109 71
rect 164 84 170 89
rect 186 89 188 91
rect 190 89 192 91
rect 164 82 166 84
rect 168 82 170 84
rect 164 81 170 82
rect 177 83 181 85
rect 177 81 178 83
rect 180 81 181 83
rect 186 84 192 89
rect 219 89 221 91
rect 223 89 225 91
rect 219 88 225 89
rect 258 89 260 91
rect 262 89 264 91
rect 258 88 264 89
rect 293 89 295 91
rect 297 89 299 91
rect 186 82 188 84
rect 190 82 192 84
rect 186 81 192 82
rect 134 77 158 81
rect 177 77 181 81
rect 223 84 243 85
rect 223 82 239 84
rect 241 82 243 84
rect 223 81 243 82
rect 293 84 299 89
rect 315 89 317 91
rect 319 89 321 91
rect 293 82 295 84
rect 297 82 299 84
rect 293 81 299 82
rect 306 83 310 85
rect 306 81 307 83
rect 309 81 310 83
rect 315 84 321 89
rect 315 82 317 84
rect 319 82 321 84
rect 315 81 321 82
rect 94 67 96 69
rect 98 67 100 69
rect 94 61 100 67
rect 132 73 138 77
rect 154 76 194 77
rect 154 74 178 76
rect 180 74 194 76
rect 81 60 100 61
rect 81 58 83 60
rect 85 58 100 60
rect 81 57 100 58
rect 78 46 79 48
rect 90 44 94 57
rect 132 63 136 73
rect 142 72 146 74
rect 154 73 194 74
rect 142 70 143 72
rect 145 70 146 72
rect 142 69 146 70
rect 132 61 133 63
rect 135 61 136 63
rect 132 59 136 61
rect 139 65 146 69
rect 139 54 143 65
rect 182 60 186 65
rect 182 58 183 60
rect 185 58 186 60
rect 125 53 143 54
rect 125 51 127 53
rect 129 52 143 53
rect 129 51 154 52
rect 125 50 150 51
rect 139 49 150 50
rect 152 49 154 51
rect 139 48 154 49
rect 159 51 163 53
rect 159 49 160 51
rect 162 49 163 51
rect 159 44 163 49
rect 182 56 186 58
rect 190 62 194 73
rect 190 60 196 62
rect 190 58 193 60
rect 195 58 196 60
rect 190 56 196 58
rect 190 53 194 56
rect 174 49 194 53
rect 174 45 178 49
rect 90 43 109 44
rect 90 41 105 43
rect 107 41 109 43
rect 90 40 109 41
rect 138 43 160 44
rect 129 40 133 42
rect 138 41 140 43
rect 142 42 160 43
rect 162 42 163 44
rect 142 41 163 42
rect 168 44 178 45
rect 168 42 170 44
rect 172 42 178 44
rect 168 41 178 42
rect 211 78 212 81
rect 223 77 227 81
rect 215 73 227 77
rect 215 61 219 73
rect 263 77 287 81
rect 306 77 310 81
rect 215 59 216 61
rect 218 59 219 61
rect 215 54 219 59
rect 261 73 267 77
rect 283 76 323 77
rect 283 74 307 76
rect 309 74 323 76
rect 261 63 265 73
rect 271 72 275 74
rect 283 73 323 74
rect 271 70 272 72
rect 274 70 275 72
rect 271 69 275 70
rect 261 61 262 63
rect 264 61 265 63
rect 261 59 265 61
rect 268 65 275 69
rect 215 50 232 54
rect 138 40 163 41
rect 129 38 130 40
rect 132 38 133 40
rect 129 35 133 38
rect 185 37 191 38
rect 185 35 187 37
rect 189 35 191 37
rect 217 46 223 47
rect 217 44 219 46
rect 221 44 223 46
rect 217 35 223 44
rect 228 46 232 50
rect 228 44 229 46
rect 231 44 232 46
rect 228 42 232 44
rect 237 46 243 47
rect 237 44 239 46
rect 241 44 243 46
rect 237 35 243 44
rect 268 54 272 65
rect 311 60 315 65
rect 311 58 312 60
rect 314 58 315 60
rect 254 53 272 54
rect 311 56 315 58
rect 319 62 323 73
rect 319 60 325 62
rect 319 58 322 60
rect 324 58 325 60
rect 319 56 325 58
rect 319 53 323 56
rect 254 51 256 53
rect 258 52 272 53
rect 258 51 283 52
rect 254 50 279 51
rect 268 49 279 50
rect 281 49 283 51
rect 268 48 283 49
rect 288 51 292 53
rect 288 49 289 51
rect 291 49 292 51
rect 288 44 292 49
rect 303 49 323 53
rect 303 45 307 49
rect 267 43 289 44
rect 258 40 262 42
rect 267 41 269 43
rect 271 42 289 43
rect 291 42 292 44
rect 271 41 292 42
rect 297 44 307 45
rect 297 42 299 44
rect 301 42 307 44
rect 297 41 307 42
rect 345 65 346 71
rect 349 70 353 91
rect 372 73 376 91
rect 395 89 397 91
rect 399 89 401 91
rect 395 88 401 89
rect 430 89 432 91
rect 434 89 436 91
rect 372 71 373 73
rect 375 71 376 73
rect 349 69 357 70
rect 349 67 353 69
rect 355 67 357 69
rect 349 66 357 67
rect 361 69 367 70
rect 372 69 376 71
rect 430 84 436 89
rect 452 89 454 91
rect 456 89 458 91
rect 430 82 432 84
rect 434 82 436 84
rect 430 81 436 82
rect 443 83 447 85
rect 443 81 444 83
rect 446 81 447 83
rect 452 84 458 89
rect 485 89 487 91
rect 489 89 491 91
rect 485 88 491 89
rect 524 89 526 91
rect 528 89 530 91
rect 524 88 530 89
rect 559 89 561 91
rect 563 89 565 91
rect 452 82 454 84
rect 456 82 458 84
rect 452 81 458 82
rect 400 77 424 81
rect 443 77 447 81
rect 489 84 509 85
rect 489 82 505 84
rect 507 82 509 84
rect 489 81 509 82
rect 559 84 565 89
rect 581 89 583 91
rect 585 89 587 91
rect 559 82 561 84
rect 563 82 565 84
rect 559 81 565 82
rect 572 83 576 85
rect 572 81 573 83
rect 575 81 576 83
rect 581 84 587 89
rect 581 82 583 84
rect 585 82 587 84
rect 581 81 587 82
rect 361 67 363 69
rect 365 67 367 69
rect 361 61 367 67
rect 398 73 404 77
rect 420 76 460 77
rect 420 74 444 76
rect 446 74 460 76
rect 348 60 367 61
rect 348 58 350 60
rect 352 58 367 60
rect 348 57 367 58
rect 345 46 346 48
rect 267 40 292 41
rect 357 44 361 57
rect 398 63 402 73
rect 408 72 412 74
rect 420 73 460 74
rect 408 70 409 72
rect 411 70 412 72
rect 408 69 412 70
rect 398 61 399 63
rect 401 61 402 63
rect 398 59 402 61
rect 405 65 412 69
rect 405 54 409 65
rect 448 60 452 65
rect 448 58 449 60
rect 451 58 452 60
rect 391 53 409 54
rect 391 51 393 53
rect 395 52 409 53
rect 395 51 420 52
rect 391 50 416 51
rect 405 49 416 50
rect 418 49 420 51
rect 405 48 420 49
rect 425 51 429 53
rect 425 49 426 51
rect 428 49 429 51
rect 425 44 429 49
rect 448 56 452 58
rect 456 62 460 73
rect 456 60 462 62
rect 456 58 459 60
rect 461 58 462 60
rect 456 56 462 58
rect 456 53 460 56
rect 440 49 460 53
rect 440 45 444 49
rect 357 43 376 44
rect 357 41 372 43
rect 374 41 376 43
rect 357 40 376 41
rect 404 43 426 44
rect 395 40 399 42
rect 404 41 406 43
rect 408 42 426 43
rect 428 42 429 44
rect 408 41 429 42
rect 434 44 444 45
rect 434 42 436 44
rect 438 42 444 44
rect 434 41 444 42
rect 477 78 478 81
rect 489 77 493 81
rect 481 73 493 77
rect 481 61 485 73
rect 529 77 553 81
rect 572 77 576 81
rect 481 59 482 61
rect 484 59 485 61
rect 481 54 485 59
rect 527 73 533 77
rect 549 76 589 77
rect 549 74 573 76
rect 575 74 589 76
rect 527 63 531 73
rect 537 72 541 74
rect 549 73 589 74
rect 537 70 538 72
rect 540 70 541 72
rect 537 69 541 70
rect 527 61 528 63
rect 530 61 531 63
rect 527 59 531 61
rect 534 65 541 69
rect 481 50 498 54
rect 404 40 429 41
rect 483 46 489 47
rect 483 44 485 46
rect 487 44 489 46
rect 258 38 259 40
rect 261 38 262 40
rect 395 38 396 40
rect 398 38 399 40
rect 258 35 262 38
rect 314 37 320 38
rect 314 35 316 37
rect 318 35 320 37
rect 395 35 399 38
rect 451 37 457 38
rect 451 35 453 37
rect 455 35 457 37
rect 483 35 489 44
rect 494 46 498 50
rect 494 44 495 46
rect 497 44 498 46
rect 494 42 498 44
rect 503 46 509 47
rect 503 44 505 46
rect 507 44 509 46
rect 503 35 509 44
rect 534 54 538 65
rect 577 60 581 65
rect 577 58 578 60
rect 580 58 581 60
rect 520 53 538 54
rect 520 51 522 53
rect 524 52 538 53
rect 524 51 549 52
rect 520 50 545 51
rect 534 49 545 50
rect 547 49 549 51
rect 534 48 549 49
rect 554 51 558 53
rect 554 49 555 51
rect 557 49 558 51
rect 554 44 558 49
rect 577 56 581 58
rect 585 62 589 73
rect 585 60 591 62
rect 585 58 588 60
rect 590 58 591 60
rect 585 56 591 58
rect 585 53 589 56
rect 569 49 589 53
rect 569 45 573 49
rect 533 43 555 44
rect 524 40 528 42
rect 533 41 535 43
rect 537 42 555 43
rect 557 42 558 44
rect 537 41 558 42
rect 563 44 573 45
rect 563 42 565 44
rect 567 42 573 44
rect 563 41 573 42
rect 612 65 613 71
rect 616 70 620 91
rect 639 73 643 91
rect 661 89 663 91
rect 665 89 667 91
rect 661 88 667 89
rect 696 89 698 91
rect 700 89 702 91
rect 639 71 640 73
rect 642 71 643 73
rect 616 69 624 70
rect 616 67 620 69
rect 622 67 624 69
rect 616 66 624 67
rect 628 69 634 70
rect 639 69 643 71
rect 696 84 702 89
rect 718 89 720 91
rect 722 89 724 91
rect 696 82 698 84
rect 700 82 702 84
rect 696 81 702 82
rect 709 83 713 85
rect 709 81 710 83
rect 712 81 713 83
rect 718 84 724 89
rect 751 89 753 91
rect 755 89 757 91
rect 751 88 757 89
rect 790 89 792 91
rect 794 89 796 91
rect 790 88 796 89
rect 825 89 827 91
rect 829 89 831 91
rect 718 82 720 84
rect 722 82 724 84
rect 718 81 724 82
rect 666 77 690 81
rect 709 77 713 81
rect 755 84 775 85
rect 755 82 771 84
rect 773 82 775 84
rect 755 81 775 82
rect 825 84 831 89
rect 847 89 849 91
rect 851 89 853 91
rect 825 82 827 84
rect 829 82 831 84
rect 825 81 831 82
rect 838 83 842 85
rect 838 81 839 83
rect 841 81 842 83
rect 847 84 853 89
rect 847 82 849 84
rect 851 82 853 84
rect 847 81 853 82
rect 628 67 630 69
rect 632 67 634 69
rect 628 61 634 67
rect 664 73 670 77
rect 686 76 726 77
rect 686 74 710 76
rect 712 74 726 76
rect 615 60 634 61
rect 615 58 617 60
rect 619 58 634 60
rect 615 57 634 58
rect 612 46 613 48
rect 533 40 558 41
rect 624 44 628 57
rect 664 63 668 73
rect 674 72 678 74
rect 686 73 726 74
rect 674 70 675 72
rect 677 70 678 72
rect 674 69 678 70
rect 664 61 665 63
rect 667 61 668 63
rect 664 59 668 61
rect 671 65 678 69
rect 671 54 675 65
rect 714 60 718 65
rect 714 58 715 60
rect 717 58 718 60
rect 657 53 675 54
rect 657 51 659 53
rect 661 52 675 53
rect 661 51 686 52
rect 657 50 682 51
rect 671 49 682 50
rect 684 49 686 51
rect 671 48 686 49
rect 691 51 695 53
rect 691 49 692 51
rect 694 49 695 51
rect 691 44 695 49
rect 714 56 718 58
rect 722 62 726 73
rect 722 60 728 62
rect 722 58 725 60
rect 727 58 728 60
rect 722 56 728 58
rect 722 53 726 56
rect 706 49 726 53
rect 706 45 710 49
rect 624 43 643 44
rect 624 41 639 43
rect 641 41 643 43
rect 624 40 643 41
rect 670 43 692 44
rect 661 40 665 42
rect 670 41 672 43
rect 674 42 692 43
rect 694 42 695 44
rect 674 41 695 42
rect 700 44 710 45
rect 700 42 702 44
rect 704 42 710 44
rect 700 41 710 42
rect 743 78 744 81
rect 755 77 759 81
rect 747 73 759 77
rect 747 61 751 73
rect 795 77 819 81
rect 838 77 842 81
rect 747 59 748 61
rect 750 59 751 61
rect 747 54 751 59
rect 793 73 799 77
rect 815 76 855 77
rect 815 74 839 76
rect 841 74 855 76
rect 793 63 797 73
rect 803 72 807 74
rect 815 73 855 74
rect 803 70 804 72
rect 806 70 807 72
rect 803 69 807 70
rect 793 61 794 63
rect 796 61 797 63
rect 793 59 797 61
rect 800 65 807 69
rect 747 50 764 54
rect 749 46 755 47
rect 749 44 751 46
rect 753 44 755 46
rect 670 40 695 41
rect 524 38 525 40
rect 527 38 528 40
rect 661 38 662 40
rect 664 38 665 40
rect 524 35 528 38
rect 580 37 586 38
rect 580 35 582 37
rect 584 35 586 37
rect 661 35 665 38
rect 717 37 723 38
rect 717 35 719 37
rect 721 35 723 37
rect 749 35 755 44
rect 760 46 764 50
rect 760 44 761 46
rect 763 44 764 46
rect 760 42 764 44
rect 769 46 775 47
rect 769 44 771 46
rect 773 44 775 46
rect 769 35 775 44
rect 800 54 804 65
rect 843 60 847 65
rect 843 58 844 60
rect 846 58 847 60
rect 786 53 804 54
rect 786 51 788 53
rect 790 52 804 53
rect 790 51 815 52
rect 786 50 811 51
rect 800 49 811 50
rect 813 49 815 51
rect 800 48 815 49
rect 820 51 824 53
rect 820 49 821 51
rect 823 49 824 51
rect 820 44 824 49
rect 843 56 847 58
rect 851 62 855 73
rect 851 60 857 62
rect 851 58 854 60
rect 856 58 857 60
rect 851 56 857 58
rect 851 53 855 56
rect 835 49 855 53
rect 835 45 839 49
rect 799 43 821 44
rect 790 40 794 42
rect 799 41 801 43
rect 803 42 821 43
rect 823 42 824 44
rect 803 41 824 42
rect 829 44 839 45
rect 829 42 831 44
rect 833 42 839 44
rect 829 41 839 42
rect 877 65 878 71
rect 881 70 885 91
rect 904 73 908 91
rect 904 71 905 73
rect 907 71 908 73
rect 881 69 889 70
rect 881 67 885 69
rect 887 67 889 69
rect 881 66 889 67
rect 893 69 899 70
rect 904 69 908 71
rect 893 67 895 69
rect 897 67 899 69
rect 893 61 899 67
rect 880 60 899 61
rect 880 58 882 60
rect 884 58 899 60
rect 880 57 899 58
rect 877 46 878 48
rect 799 40 824 41
rect 889 44 893 57
rect 889 43 908 44
rect 889 41 904 43
rect 906 41 908 43
rect 889 40 908 41
rect 790 38 791 40
rect 793 38 794 40
rect 790 35 794 38
rect 846 37 852 38
rect 846 35 848 37
rect 850 35 852 37
<< via1 >>
rect 176 364 178 366
rect 76 341 78 343
rect 104 340 106 342
rect 124 331 126 333
rect 407 364 409 366
rect 234 348 236 350
rect 162 323 164 325
rect 255 349 257 351
rect 224 331 226 333
rect 265 340 267 342
rect 280 348 282 350
rect 297 349 299 351
rect 305 340 307 342
rect 333 340 335 342
rect 384 349 386 351
rect 353 332 355 334
rect 458 348 460 350
rect 479 349 481 351
rect 448 331 450 333
rect 489 340 491 342
rect 504 348 506 350
rect 521 349 523 351
rect 529 340 531 342
rect 561 340 563 342
rect 608 349 610 351
rect 577 331 579 333
rect 656 339 658 341
rect 705 352 707 354
rect 673 333 675 335
rect 742 364 744 366
rect 724 334 726 336
rect 791 364 793 366
rect 773 336 775 338
rect 841 364 843 366
rect 823 335 825 337
rect 94 270 96 272
rect 76 243 78 245
rect 144 270 146 272
rect 126 245 128 247
rect 344 270 346 272
rect 326 242 328 244
rect 394 270 396 272
rect 376 245 378 247
rect 438 270 440 272
rect 494 270 496 272
rect 476 239 478 241
rect 544 270 546 272
rect 526 241 528 243
rect 594 270 596 272
rect 576 242 578 244
rect 650 270 652 272
rect 626 244 628 246
rect 701 246 703 248
rect 717 246 719 248
rect 749 230 751 232
rect 801 246 803 248
rect 818 237 820 239
rect 76 155 78 157
rect 155 161 157 163
rect 124 143 126 145
rect 165 169 167 171
rect 180 160 182 162
rect 197 161 199 163
rect 205 152 207 154
rect 233 152 235 154
rect 284 161 286 163
rect 253 146 255 148
rect 300 141 302 143
rect 379 161 381 163
rect 348 143 350 145
rect 404 160 406 162
rect 421 161 423 163
rect 429 152 431 154
rect 457 152 459 154
rect 508 161 510 163
rect 477 146 479 148
rect 603 161 605 163
rect 572 143 574 145
rect 525 136 527 138
rect 628 160 630 162
rect 645 161 647 163
rect 653 152 655 154
rect 681 152 683 154
rect 732 161 734 163
rect 701 144 703 146
rect 766 176 768 178
rect 748 144 750 146
rect 147 58 149 60
rect 198 67 200 69
rect 167 49 169 51
rect 223 66 225 68
rect 240 67 242 69
rect 248 58 250 60
rect 198 29 200 31
rect 276 58 278 60
rect 327 67 329 69
rect 296 51 298 53
rect 360 82 362 84
rect 342 51 344 53
rect 413 58 415 60
rect 464 67 466 69
rect 433 49 435 51
rect 489 66 491 68
rect 506 67 508 69
rect 514 58 516 60
rect 219 29 221 31
rect 461 29 463 31
rect 542 58 544 60
rect 593 67 595 69
rect 562 50 564 52
rect 627 82 629 84
rect 609 50 611 52
rect 708 66 710 68
rect 730 67 732 69
rect 699 49 701 51
rect 755 66 757 68
rect 772 67 774 69
rect 780 58 782 60
rect 487 29 489 31
rect 729 29 731 31
rect 808 58 810 60
rect 859 67 861 69
rect 828 49 830 51
rect 892 82 894 84
rect 874 50 876 52
rect 757 30 759 32
rect 740 14 742 16
rect 473 10 475 12
<< via2 >>
rect 743 382 745 384
rect 792 382 794 384
rect 842 382 844 384
rect 271 301 273 303
rect 94 288 96 290
rect 144 288 146 290
rect 121 245 123 247
rect 344 275 346 277
rect 439 289 441 291
rect 400 270 402 272
rect 500 270 502 272
rect 512 270 514 272
rect 529 270 531 272
rect 600 270 602 272
rect 630 270 632 272
rect 76 207 78 209
rect 476 210 478 212
rect 718 210 720 212
rect 750 210 752 212
rect 291 199 293 201
rect 165 195 167 197
rect 358 195 360 197
rect 441 195 443 197
rect 517 195 519 197
rect 234 130 236 132
rect 582 196 584 198
rect 817 203 819 205
rect 639 197 641 199
rect 871 203 873 205
rect 830 176 832 178
rect 300 117 302 119
rect 525 102 527 104
rect 790 100 792 102
rect 893 101 895 103
rect 345 82 347 84
rect 610 82 612 84
rect 277 20 279 22
rect 146 -6 148 -4
rect 543 18 545 20
rect 450 10 452 12
rect 500 11 502 13
rect 631 10 633 12
rect 808 -20 810 -18
<< via3 >>
rect 335 382 337 384
rect 601 210 603 212
rect 337 82 339 84
rect 601 82 603 84
<< labels >>
rlabel alu1 121 313 121 313 6 vss
rlabel alu1 177 341 177 341 6 so
rlabel alu1 221 313 221 313 6 vss
rlabel alu1 221 377 221 377 6 vdd
rlabel alu1 233 349 233 349 1 ci
rlabel alu1 93 283 93 283 6 vdd
rlabel alu1 93 219 93 219 6 vss
rlabel alu1 143 219 143 219 6 vss
rlabel alu1 143 283 143 283 6 vdd
rlabel alu1 343 219 343 219 6 vss
rlabel alu1 343 283 343 283 6 vdd
rlabel alu1 393 219 393 219 6 vss
rlabel alu1 393 283 393 283 6 vdd
rlabel alu1 493 219 493 219 6 vss
rlabel alu1 493 283 493 283 6 vdd
rlabel alu1 543 219 543 219 6 vss
rlabel alu1 543 283 543 283 6 vdd
rlabel alu1 593 219 593 219 6 vss
rlabel alu1 593 283 593 283 6 vdd
rlabel alu1 643 219 643 219 6 vss
rlabel alu1 643 283 643 283 6 vdd
rlabel alu1 445 377 445 377 6 vdd
rlabel alu1 670 377 670 377 6 vdd
rlabel alu1 254 149 254 149 6 a
rlabel alu1 246 161 246 161 6 b
rlabel alu1 121 189 121 189 6 vdd
rlabel alu1 121 125 121 125 6 vss
rlabel alu1 478 149 478 149 6 a
rlabel alu1 470 161 470 161 6 b
rlabel alu1 345 189 345 189 6 vdd
rlabel alu1 345 125 345 125 6 vss
rlabel alu1 569 189 569 189 6 vdd
rlabel alu1 569 125 569 125 6 vss
rlabel alu1 715 219 715 219 6 vss
rlabel alu1 715 283 715 283 6 vdd
rlabel alu1 92 31 92 31 6 vss
rlabel alu1 92 95 92 95 6 vdd
rlabel alu1 164 95 164 95 6 vdd
rlabel alu1 164 31 164 31 6 vss
rlabel alu1 359 31 359 31 6 vss
rlabel alu1 359 95 359 95 6 vdd
rlabel alu1 430 31 430 31 6 vss
rlabel alu1 430 95 430 95 6 vdd
rlabel alu1 626 31 626 31 6 vss
rlabel alu1 626 95 626 95 6 vdd
rlabel alu1 741 59 741 59 1 co
rlabel alu1 829 55 829 55 6 a
rlabel alu1 821 67 821 67 6 b
rlabel alu1 696 95 696 95 6 vdd
rlabel alu1 696 31 696 31 6 vss
rlabel alu1 765 125 765 125 6 vss
rlabel alu1 765 189 765 189 6 vdd
rlabel alu1 815 219 815 219 6 vss
rlabel alu1 815 283 815 283 6 vdd
rlabel alu1 741 313 741 313 6 vss
rlabel alu1 741 377 741 377 6 vdd
rlabel alu1 891 31 891 31 6 vss
rlabel alu1 891 95 891 95 6 vdd
rlabel alu1 790 313 790 313 6 vss
rlabel alu1 790 377 790 377 6 vdd
rlabel alu1 840 313 840 313 6 vss
rlabel alu1 840 377 840 377 6 vdd
rlabel polyct1 95 271 95 271 1 x3
rlabel polyct1 104 239 104 239 1 y1
rlabel alu1 77 248 77 248 1 x3y1
rlabel polyct1 354 239 354 239 1 y0
rlabel polyct1 345 271 345 271 1 x3
rlabel polyct1 395 271 395 271 1 x2
rlabel polyct1 404 239 404 239 1 y1
rlabel alu1 327 249 327 249 1 x3y0
rlabel alu1 377 250 377 250 1 x2y1
rlabel polyct1 545 271 545 271 1 x2
rlabel polyct1 554 239 554 239 1 y0
rlabel polyct1 595 271 595 271 1 x1
rlabel polyct1 604 239 604 239 1 y1
rlabel polyct1 645 271 645 271 1 x1
rlabel polyct1 654 239 654 239 1 y0
rlabel polyct1 743 365 743 365 1 x0
rlabel polyct1 752 333 752 333 1 y1
rlabel polyct1 145 271 145 271 1 x3
rlabel polyct1 154 239 154 239 1 y2
rlabel polyct1 495 271 495 271 1 x2
rlabel polyct1 504 239 504 239 1 y2
rlabel polyct1 776 145 776 145 1 y2
rlabel polyct1 767 177 767 177 1 x1
rlabel polyct1 842 365 842 365 1 x0
rlabel polyct1 851 333 851 333 1 y2
rlabel polyct1 792 365 792 365 1 x0
rlabel polyct1 801 333 801 333 1 y3
rlabel polyct1 361 83 361 83 1 x3
rlabel polyct1 370 51 370 51 1 y3
rlabel polyct1 628 83 628 83 1 x2
rlabel polyct1 637 51 637 51 1 y3
rlabel polyct1 893 83 893 83 1 x1
rlabel polyct1 902 51 902 51 1 y3
rlabel alu1 626 332 626 332 1 z1
rlabel alu1 771 241 771 241 1 z2
rlabel alu1 671 240 671 240 1 z3
rlabel alu1 652 52 652 52 1 z4
rlabel alu1 386 52 386 52 1 z5
rlabel alu1 120 51 120 51 1 z6
rlabel alu1 209 35 209 35 1 z7
rlabel alu1 121 377 121 377 6 vdd
rlabel alu1 214 220 214 220 6 vss
rlabel alu1 214 284 214 284 6 vdd
rlabel alu1 255 284 255 284 6 vdd
rlabel alu1 255 220 255 220 6 vss
rlabel alu1 437 219 437 219 6 vss
rlabel alu1 437 283 437 283 6 vdd
rlabel polyct1 439 271 439 271 1 x0
rlabel polyct1 448 239 448 239 1 y0
rlabel alu1 725 340 725 340 1 z0
<< end >>
