magic
tech scmos
timestamp 1636287559
<< ab >>
rect 265 127 305 199
rect 308 186 348 199
rect 308 182 333 186
rect 317 180 333 182
rect 338 180 348 186
rect 317 178 348 180
rect 308 127 348 178
rect 351 186 391 199
rect 351 178 368 186
rect 381 180 391 186
rect 376 178 391 180
rect 351 127 391 178
rect 394 127 434 199
rect 264 53 356 103
rect 264 31 351 53
rect 355 31 356 53
rect 358 31 456 103
rect -255 -115 -215 -43
rect -212 -56 -172 -43
rect -212 -60 -187 -56
rect -203 -62 -187 -60
rect -182 -62 -172 -56
rect -203 -64 -172 -62
rect -212 -115 -172 -64
rect -169 -56 -129 -43
rect -169 -64 -152 -56
rect -139 -62 -129 -56
rect -144 -64 -129 -62
rect -169 -115 -129 -64
rect -126 -115 -86 -43
rect 14 -127 101 -84
rect 14 -130 55 -127
rect 59 -130 101 -127
rect -256 -211 -164 -139
rect -162 -211 -64 -139
rect 14 -156 101 -130
rect 105 -122 232 -84
rect 105 -131 142 -122
rect 145 -131 232 -122
rect 105 -135 232 -131
rect 105 -137 143 -135
rect 145 -137 232 -135
rect 105 -156 232 -137
rect 234 -122 361 -84
rect 234 -131 321 -122
rect 324 -131 361 -122
rect 234 -135 361 -131
rect 234 -137 321 -135
rect 323 -137 361 -135
rect 234 -156 361 -137
rect 365 -156 539 -84
rect 543 -114 765 -84
rect 543 -122 712 -114
rect 543 -131 580 -122
rect 583 -131 712 -122
rect 543 -135 712 -131
rect 543 -137 581 -135
rect 583 -137 712 -135
rect 543 -156 712 -137
rect 716 -156 765 -114
rect 398 -290 438 -218
rect 441 -231 481 -218
rect 441 -235 466 -231
rect 450 -237 466 -235
rect 471 -237 481 -231
rect 450 -239 481 -237
rect 441 -290 481 -239
rect 484 -231 524 -218
rect 484 -239 501 -231
rect 514 -237 524 -231
rect 509 -239 524 -237
rect 484 -290 524 -239
rect 527 -290 567 -218
rect -254 -367 -214 -295
rect -211 -308 -171 -295
rect -211 -312 -186 -308
rect -202 -314 -186 -312
rect -181 -314 -171 -308
rect -202 -316 -171 -314
rect -211 -367 -171 -316
rect -168 -308 -128 -295
rect -168 -316 -151 -308
rect -138 -314 -128 -308
rect -143 -316 -128 -314
rect -168 -367 -128 -316
rect -125 -367 -85 -295
rect 397 -386 489 -314
rect 491 -386 589 -314
rect -255 -457 -163 -391
rect -255 -462 -247 -457
rect -233 -462 -163 -457
rect -255 -463 -163 -462
rect -161 -463 -63 -391
rect 16 -541 103 -469
rect 107 -507 234 -469
rect 107 -516 144 -507
rect 147 -516 234 -507
rect 107 -520 234 -516
rect 107 -522 145 -520
rect 147 -522 234 -520
rect 107 -541 234 -522
rect 236 -507 363 -469
rect 236 -516 323 -507
rect 326 -516 363 -507
rect 236 -520 363 -516
rect 236 -522 323 -520
rect 325 -522 363 -520
rect 236 -541 363 -522
rect 367 -541 541 -469
rect 545 -507 767 -469
rect 545 -516 582 -507
rect 585 -516 767 -507
rect 545 -520 767 -516
rect 545 -522 583 -520
rect 585 -522 767 -520
rect 545 -541 767 -522
rect -251 -675 -164 -603
rect -160 -641 -33 -603
rect -160 -650 -123 -641
rect -120 -650 -33 -641
rect -160 -654 -33 -650
rect -160 -656 -122 -654
rect -120 -656 -33 -654
rect -160 -675 -33 -656
rect -31 -641 96 -603
rect -31 -650 56 -641
rect 59 -650 96 -641
rect -31 -654 96 -650
rect -31 -656 56 -654
rect 58 -656 96 -654
rect -31 -675 96 -656
rect 100 -675 274 -603
rect 278 -641 500 -603
rect 278 -650 315 -641
rect 318 -650 500 -641
rect 278 -654 500 -650
rect 278 -656 316 -654
rect 318 -656 500 -654
rect 278 -675 500 -656
<< nwell >>
rect 263 159 436 204
rect 262 63 456 108
rect -257 -83 -84 -38
rect 14 -124 765 -79
rect -258 -179 -64 -134
rect 396 -258 569 -213
rect -256 -335 -83 -290
rect 395 -354 589 -309
rect -257 -431 -63 -386
rect 16 -509 767 -464
rect -251 -643 500 -598
<< pwell >>
rect 263 122 436 159
rect 262 26 456 63
rect -257 -120 -84 -83
rect 14 -161 765 -124
rect -258 -216 -64 -179
rect 396 -295 569 -258
rect -256 -372 -83 -335
rect 395 -391 589 -354
rect -257 -468 -63 -431
rect 16 -546 767 -509
rect -251 -680 500 -643
<< poly >>
rect 305 202 850 204
rect 305 188 307 202
rect -43 186 286 188
rect 305 186 331 188
rect 337 186 417 188
rect -43 185 236 186
rect -267 -41 -212 -38
rect -267 -281 -265 -41
rect -215 -54 -212 -41
rect -215 -56 -189 -54
rect -183 -56 -103 -54
rect -236 -58 -230 -56
rect -236 -60 -234 -58
rect -232 -60 -230 -58
rect -246 -65 -244 -60
rect -236 -62 -230 -60
rect -215 -62 -213 -56
rect -193 -58 -187 -56
rect -193 -60 -191 -58
rect -189 -60 -187 -58
rect -236 -67 -234 -62
rect -226 -64 -213 -62
rect -226 -67 -224 -64
rect -203 -65 -201 -60
rect -193 -62 -187 -60
rect -193 -67 -191 -62
rect -183 -67 -181 -56
rect -107 -58 -101 -56
rect -107 -60 -105 -58
rect -103 -60 -101 -58
rect -160 -65 -158 -60
rect -150 -67 -148 -63
rect -140 -67 -138 -62
rect -117 -65 -115 -60
rect -107 -62 -101 -60
rect -107 -67 -105 -62
rect -97 -67 -95 -62
rect -246 -80 -244 -77
rect -236 -80 -234 -77
rect -246 -82 -240 -80
rect -246 -84 -244 -82
rect -242 -84 -240 -82
rect -236 -83 -232 -80
rect -246 -86 -240 -84
rect -246 -94 -244 -86
rect -234 -97 -232 -83
rect -226 -88 -224 -77
rect -203 -80 -201 -77
rect -193 -80 -191 -77
rect -203 -82 -197 -80
rect -203 -84 -201 -82
rect -199 -84 -197 -82
rect -193 -83 -189 -80
rect -203 -86 -197 -84
rect -227 -90 -221 -88
rect -227 -92 -225 -90
rect -223 -92 -221 -90
rect -227 -94 -221 -92
rect -203 -94 -201 -86
rect -227 -97 -225 -94
rect -246 -104 -244 -100
rect -191 -97 -189 -83
rect -183 -88 -181 -77
rect -160 -80 -158 -77
rect -150 -80 -148 -77
rect -160 -82 -154 -80
rect -160 -84 -158 -82
rect -156 -84 -154 -82
rect -150 -83 -146 -80
rect -160 -86 -154 -84
rect -184 -90 -178 -88
rect -184 -92 -182 -90
rect -180 -92 -178 -90
rect -184 -94 -178 -92
rect -160 -94 -158 -86
rect -184 -97 -182 -94
rect -203 -104 -201 -100
rect -148 -97 -146 -83
rect -140 -88 -138 -77
rect -117 -80 -115 -77
rect -107 -80 -105 -77
rect -117 -82 -111 -80
rect -117 -84 -115 -82
rect -113 -84 -111 -82
rect -107 -83 -103 -80
rect -117 -86 -111 -84
rect -141 -90 -135 -88
rect -141 -92 -139 -90
rect -137 -92 -135 -90
rect -141 -94 -135 -92
rect -117 -94 -115 -86
rect -141 -97 -139 -94
rect -160 -104 -158 -100
rect -105 -97 -103 -83
rect -97 -88 -95 -77
rect -98 -90 -92 -88
rect -98 -92 -96 -90
rect -94 -92 -92 -90
rect -98 -94 -92 -92
rect -98 -97 -96 -94
rect -117 -104 -115 -100
rect -234 -118 -232 -106
rect -227 -111 -225 -106
rect -191 -111 -189 -106
rect -184 -111 -182 -106
rect -148 -118 -146 -106
rect -141 -118 -139 -106
rect -105 -111 -103 -106
rect -98 -118 -96 -106
rect -234 -120 -145 -118
rect -141 -120 -52 -118
rect -247 -145 -245 -141
rect -224 -148 -222 -143
rect -217 -148 -215 -143
rect -199 -145 -197 -141
rect -189 -145 -187 -141
rect -179 -145 -177 -141
rect -145 -145 -143 -141
rect -135 -145 -133 -141
rect -125 -145 -123 -141
rect -234 -157 -232 -152
rect -247 -183 -245 -170
rect -234 -173 -232 -170
rect -107 -148 -105 -143
rect -100 -148 -98 -143
rect -77 -145 -75 -141
rect -90 -157 -88 -152
rect -90 -173 -88 -170
rect -241 -175 -232 -173
rect -241 -177 -239 -175
rect -237 -177 -235 -175
rect -224 -176 -222 -173
rect -217 -176 -215 -173
rect -199 -176 -197 -173
rect -189 -176 -187 -173
rect -179 -176 -177 -173
rect -145 -176 -143 -173
rect -135 -176 -133 -173
rect -125 -176 -123 -173
rect -107 -176 -105 -173
rect -100 -176 -98 -173
rect -90 -175 -81 -173
rect -241 -179 -235 -177
rect -247 -185 -241 -183
rect -247 -187 -245 -185
rect -243 -187 -241 -185
rect -247 -189 -241 -187
rect -247 -192 -245 -189
rect -237 -192 -235 -179
rect -227 -178 -221 -176
rect -227 -180 -225 -178
rect -223 -180 -221 -178
rect -227 -182 -221 -180
rect -217 -178 -195 -176
rect -217 -180 -206 -178
rect -204 -180 -199 -178
rect -197 -180 -195 -178
rect -217 -182 -195 -180
rect -191 -178 -185 -176
rect -191 -180 -189 -178
rect -187 -180 -185 -178
rect -191 -182 -185 -180
rect -181 -178 -175 -176
rect -181 -180 -179 -178
rect -177 -180 -175 -178
rect -181 -182 -175 -180
rect -147 -178 -141 -176
rect -147 -180 -145 -178
rect -143 -180 -141 -178
rect -147 -182 -141 -180
rect -137 -178 -131 -176
rect -137 -180 -135 -178
rect -133 -180 -131 -178
rect -137 -182 -131 -180
rect -127 -178 -105 -176
rect -127 -180 -125 -178
rect -123 -180 -118 -178
rect -116 -180 -105 -178
rect -127 -182 -105 -180
rect -101 -178 -95 -176
rect -101 -180 -99 -178
rect -97 -180 -95 -178
rect -101 -182 -95 -180
rect -227 -185 -225 -182
rect -217 -185 -215 -182
rect -197 -185 -195 -182
rect -190 -185 -188 -182
rect -247 -209 -245 -205
rect -237 -207 -235 -202
rect -227 -204 -225 -199
rect -217 -204 -215 -199
rect -179 -191 -177 -182
rect -145 -191 -143 -182
rect -134 -185 -132 -182
rect -127 -185 -125 -182
rect -107 -185 -105 -182
rect -97 -185 -95 -182
rect -87 -177 -85 -175
rect -83 -177 -81 -175
rect -87 -179 -81 -177
rect -87 -192 -85 -179
rect -77 -183 -75 -170
rect -81 -185 -75 -183
rect -81 -187 -79 -185
rect -77 -187 -75 -185
rect -81 -189 -75 -187
rect -77 -192 -75 -189
rect -107 -204 -105 -199
rect -97 -204 -95 -199
rect -197 -209 -195 -205
rect -190 -209 -188 -205
rect -179 -209 -177 -205
rect -145 -209 -143 -205
rect -134 -209 -132 -205
rect -127 -209 -125 -205
rect -87 -207 -85 -202
rect -77 -209 -75 -205
rect -268 -283 -210 -281
rect -212 -306 -210 -283
rect -214 -308 -188 -306
rect -182 -308 -102 -306
rect -235 -310 -229 -308
rect -235 -312 -233 -310
rect -231 -312 -229 -310
rect -245 -317 -243 -312
rect -235 -314 -229 -312
rect -214 -314 -212 -308
rect -192 -310 -186 -308
rect -192 -312 -190 -310
rect -188 -312 -186 -310
rect -235 -319 -233 -314
rect -225 -316 -212 -314
rect -225 -319 -223 -316
rect -202 -317 -200 -312
rect -192 -314 -186 -312
rect -192 -319 -190 -314
rect -182 -319 -180 -308
rect -106 -310 -100 -308
rect -106 -312 -104 -310
rect -102 -312 -100 -310
rect -159 -317 -157 -312
rect -149 -319 -147 -315
rect -139 -319 -137 -314
rect -116 -317 -114 -312
rect -106 -314 -100 -312
rect -54 -314 -52 -120
rect -106 -319 -104 -314
rect -96 -317 -52 -314
rect -96 -319 -94 -317
rect -245 -332 -243 -329
rect -235 -332 -233 -329
rect -245 -334 -239 -332
rect -245 -336 -243 -334
rect -241 -336 -239 -334
rect -235 -335 -231 -332
rect -245 -338 -239 -336
rect -245 -346 -243 -338
rect -233 -349 -231 -335
rect -225 -340 -223 -329
rect -202 -332 -200 -329
rect -192 -332 -190 -329
rect -202 -334 -196 -332
rect -202 -336 -200 -334
rect -198 -336 -196 -334
rect -192 -335 -188 -332
rect -202 -338 -196 -336
rect -226 -342 -220 -340
rect -226 -344 -224 -342
rect -222 -344 -220 -342
rect -226 -346 -220 -344
rect -202 -346 -200 -338
rect -226 -349 -224 -346
rect -245 -356 -243 -352
rect -190 -349 -188 -335
rect -182 -340 -180 -329
rect -159 -332 -157 -329
rect -149 -332 -147 -329
rect -159 -334 -153 -332
rect -159 -336 -157 -334
rect -155 -336 -153 -334
rect -149 -335 -145 -332
rect -159 -338 -153 -336
rect -183 -342 -177 -340
rect -183 -344 -181 -342
rect -179 -344 -177 -342
rect -183 -346 -177 -344
rect -159 -346 -157 -338
rect -183 -349 -181 -346
rect -202 -356 -200 -352
rect -147 -349 -145 -335
rect -139 -340 -137 -329
rect -116 -332 -114 -329
rect -106 -332 -104 -329
rect -116 -334 -110 -332
rect -116 -336 -114 -334
rect -112 -336 -110 -334
rect -106 -335 -102 -332
rect -116 -338 -110 -336
rect -140 -342 -134 -340
rect -140 -344 -138 -342
rect -136 -344 -134 -342
rect -140 -346 -134 -344
rect -116 -346 -114 -338
rect -140 -349 -138 -346
rect -159 -356 -157 -352
rect -104 -349 -102 -335
rect -96 -340 -94 -329
rect -97 -342 -91 -340
rect -97 -344 -95 -342
rect -93 -344 -91 -342
rect -97 -346 -91 -344
rect -97 -349 -95 -346
rect -116 -356 -114 -352
rect -233 -370 -231 -358
rect -226 -363 -224 -358
rect -190 -363 -188 -358
rect -183 -363 -181 -358
rect -147 -370 -145 -358
rect -140 -370 -138 -358
rect -104 -363 -102 -358
rect -97 -370 -95 -358
rect -233 -372 -144 -370
rect -140 -372 -95 -370
rect -146 -377 -144 -372
rect -43 -377 -40 185
rect 284 184 290 186
rect 284 182 286 184
rect 288 182 290 184
rect 274 177 276 182
rect 284 180 290 182
rect 305 180 307 186
rect 327 184 333 186
rect 327 182 329 184
rect 331 182 333 184
rect 284 175 286 180
rect 294 178 307 180
rect 294 175 296 178
rect 317 177 319 182
rect 327 180 333 182
rect 327 175 329 180
rect 337 175 339 186
rect 413 184 419 186
rect 413 182 415 184
rect 417 182 419 184
rect 360 177 362 182
rect 370 175 372 179
rect 380 175 382 180
rect 403 177 405 182
rect 413 180 419 182
rect 413 175 415 180
rect 423 178 830 180
rect 423 175 425 178
rect 274 162 276 165
rect 284 162 286 165
rect 274 160 280 162
rect 274 158 276 160
rect 278 158 280 160
rect 284 159 288 162
rect 274 156 280 158
rect 274 148 276 156
rect 286 145 288 159
rect 294 154 296 165
rect 317 162 319 165
rect 327 162 329 165
rect 317 160 323 162
rect 317 158 319 160
rect 321 158 323 160
rect 327 159 331 162
rect 317 156 323 158
rect 293 152 299 154
rect 293 150 295 152
rect 297 150 299 152
rect 293 148 299 150
rect 317 148 319 156
rect 293 145 295 148
rect 274 138 276 142
rect 329 145 331 159
rect 337 154 339 165
rect 360 162 362 165
rect 370 162 372 165
rect 360 160 366 162
rect 360 158 362 160
rect 364 158 366 160
rect 370 159 374 162
rect 360 156 366 158
rect 336 152 342 154
rect 336 150 338 152
rect 340 150 342 152
rect 336 148 342 150
rect 360 148 362 156
rect 336 145 338 148
rect 317 138 319 142
rect 372 145 374 159
rect 380 154 382 165
rect 403 162 405 165
rect 413 162 415 165
rect 403 160 409 162
rect 403 158 405 160
rect 407 158 409 160
rect 413 159 417 162
rect 403 156 409 158
rect 379 152 385 154
rect 379 150 381 152
rect 383 150 385 152
rect 379 148 385 150
rect 403 148 405 156
rect 379 145 381 148
rect 360 138 362 142
rect 415 145 417 159
rect 423 154 425 165
rect 422 152 428 154
rect 422 150 424 152
rect 426 150 428 152
rect 422 148 428 150
rect 422 145 424 148
rect 403 138 405 142
rect 286 124 288 136
rect 293 131 295 136
rect 329 131 331 136
rect 336 131 338 136
rect 372 124 374 136
rect 379 124 381 136
rect 415 131 417 136
rect 422 124 424 136
rect 286 122 375 124
rect 379 122 424 124
rect 273 97 275 101
rect 296 94 298 99
rect 303 94 305 99
rect 321 97 323 101
rect 331 97 333 101
rect 341 97 343 101
rect 375 97 377 101
rect 385 97 387 101
rect 395 97 397 101
rect 286 85 288 90
rect 273 59 275 72
rect 286 69 288 72
rect 413 94 415 99
rect 420 94 422 99
rect 443 97 445 101
rect 430 85 432 90
rect 430 69 432 72
rect 279 67 288 69
rect 279 65 281 67
rect 283 65 285 67
rect 296 66 298 69
rect 303 66 305 69
rect 321 66 323 69
rect 331 66 333 69
rect 341 66 343 69
rect 375 66 377 69
rect 385 66 387 69
rect 395 66 397 69
rect 413 66 415 69
rect 420 66 422 69
rect 430 67 439 69
rect 279 63 285 65
rect 273 57 279 59
rect 273 55 275 57
rect 277 55 279 57
rect 273 53 279 55
rect 273 50 275 53
rect 283 50 285 63
rect 293 64 299 66
rect 293 62 295 64
rect 297 62 299 64
rect 293 60 299 62
rect 303 64 325 66
rect 303 62 314 64
rect 316 62 321 64
rect 323 62 325 64
rect 303 60 325 62
rect 329 64 335 66
rect 329 62 331 64
rect 333 62 335 64
rect 329 60 335 62
rect 339 64 345 66
rect 339 62 341 64
rect 343 62 345 64
rect 339 60 345 62
rect 373 64 379 66
rect 373 62 375 64
rect 377 62 379 64
rect 373 60 379 62
rect 383 64 389 66
rect 383 62 385 64
rect 387 62 389 64
rect 383 60 389 62
rect 393 64 415 66
rect 393 62 395 64
rect 397 62 402 64
rect 404 62 415 64
rect 393 60 415 62
rect 419 64 425 66
rect 419 62 421 64
rect 423 62 425 64
rect 419 60 425 62
rect 293 57 295 60
rect 303 57 305 60
rect 323 57 325 60
rect 330 57 332 60
rect 273 33 275 37
rect 283 35 285 40
rect 293 38 295 43
rect 303 38 305 43
rect 341 51 343 60
rect 375 51 377 60
rect 386 57 388 60
rect 393 57 395 60
rect 413 57 415 60
rect 423 57 425 60
rect 433 65 435 67
rect 437 65 439 67
rect 433 63 439 65
rect 433 50 435 63
rect 443 59 445 72
rect 439 57 445 59
rect 439 55 441 57
rect 443 55 445 57
rect 439 53 445 55
rect 443 50 445 53
rect 413 38 415 43
rect 423 38 425 43
rect 323 33 325 37
rect 330 33 332 37
rect 341 33 343 37
rect 375 33 377 37
rect 386 33 388 37
rect 393 33 395 37
rect 433 35 435 40
rect 443 33 445 37
rect 24 -90 26 -86
rect 34 -90 36 -86
rect 44 -90 46 -86
rect 62 -93 64 -88
rect 69 -93 71 -88
rect 92 -90 94 -86
rect 112 -90 114 -86
rect 119 -90 121 -86
rect 79 -102 81 -97
rect 153 -90 155 -86
rect 163 -90 165 -86
rect 173 -90 175 -86
rect 132 -99 134 -95
rect 79 -118 81 -115
rect 24 -121 26 -118
rect 34 -121 36 -118
rect 44 -121 46 -118
rect 62 -121 64 -118
rect 69 -121 71 -118
rect 79 -120 88 -118
rect 22 -123 28 -121
rect 22 -125 24 -123
rect 26 -125 28 -123
rect 22 -127 28 -125
rect 32 -123 38 -121
rect 32 -125 34 -123
rect 36 -125 38 -123
rect 32 -127 38 -125
rect 42 -123 64 -121
rect 42 -125 44 -123
rect 46 -125 51 -123
rect 53 -125 64 -123
rect 42 -127 64 -125
rect 68 -123 74 -121
rect 68 -125 70 -123
rect 72 -125 74 -123
rect 68 -127 74 -125
rect 24 -136 26 -127
rect 35 -130 37 -127
rect 42 -130 44 -127
rect 62 -130 64 -127
rect 72 -130 74 -127
rect 82 -122 84 -120
rect 86 -122 88 -120
rect 82 -124 88 -122
rect 82 -137 84 -124
rect 92 -128 94 -115
rect 112 -121 114 -108
rect 119 -113 121 -108
rect 118 -115 124 -113
rect 118 -117 120 -115
rect 122 -117 124 -115
rect 118 -119 124 -117
rect 108 -123 114 -121
rect 108 -125 110 -123
rect 112 -125 114 -123
rect 108 -127 114 -125
rect 88 -130 94 -128
rect 88 -132 90 -130
rect 92 -132 94 -130
rect 88 -134 94 -132
rect 92 -137 94 -134
rect 112 -135 114 -127
rect 122 -135 124 -119
rect 132 -120 134 -111
rect 191 -93 193 -88
rect 198 -93 200 -88
rect 221 -90 223 -86
rect 243 -90 245 -86
rect 208 -102 210 -97
rect 266 -93 268 -88
rect 273 -93 275 -88
rect 291 -90 293 -86
rect 301 -90 303 -86
rect 311 -90 313 -86
rect 256 -102 258 -97
rect 208 -118 210 -115
rect 128 -122 134 -120
rect 153 -121 155 -118
rect 163 -121 165 -118
rect 173 -121 175 -118
rect 191 -121 193 -118
rect 198 -121 200 -118
rect 208 -120 217 -118
rect 128 -124 130 -122
rect 132 -124 134 -122
rect 128 -126 134 -124
rect 132 -135 134 -126
rect 151 -123 157 -121
rect 151 -125 153 -123
rect 155 -125 157 -123
rect 151 -127 157 -125
rect 161 -123 167 -121
rect 161 -125 163 -123
rect 165 -125 167 -123
rect 161 -127 167 -125
rect 171 -123 193 -121
rect 171 -125 173 -123
rect 175 -125 180 -123
rect 182 -125 193 -123
rect 171 -127 193 -125
rect 197 -123 203 -121
rect 197 -125 199 -123
rect 201 -125 203 -123
rect 197 -127 203 -125
rect 62 -149 64 -144
rect 72 -149 74 -144
rect 24 -154 26 -150
rect 35 -154 37 -150
rect 42 -154 44 -150
rect 82 -152 84 -147
rect 153 -136 155 -127
rect 164 -130 166 -127
rect 171 -130 173 -127
rect 191 -130 193 -127
rect 201 -130 203 -127
rect 211 -122 213 -120
rect 215 -122 217 -120
rect 211 -124 217 -122
rect 112 -145 114 -141
rect 122 -145 124 -141
rect 132 -145 134 -141
rect 92 -154 94 -150
rect 211 -137 213 -124
rect 221 -128 223 -115
rect 217 -130 223 -128
rect 217 -132 219 -130
rect 221 -132 223 -130
rect 217 -134 223 -132
rect 221 -137 223 -134
rect 243 -128 245 -115
rect 256 -118 258 -115
rect 345 -90 347 -86
rect 352 -90 354 -86
rect 372 -90 374 -86
rect 332 -99 334 -95
rect 249 -120 258 -118
rect 249 -122 251 -120
rect 253 -122 255 -120
rect 266 -121 268 -118
rect 273 -121 275 -118
rect 291 -121 293 -118
rect 301 -121 303 -118
rect 311 -121 313 -118
rect 332 -120 334 -111
rect 345 -113 347 -108
rect 342 -115 348 -113
rect 342 -117 344 -115
rect 346 -117 348 -115
rect 342 -119 348 -117
rect 249 -124 255 -122
rect 243 -130 249 -128
rect 243 -132 245 -130
rect 247 -132 249 -130
rect 243 -134 249 -132
rect 243 -137 245 -134
rect 253 -137 255 -124
rect 263 -123 269 -121
rect 263 -125 265 -123
rect 267 -125 269 -123
rect 263 -127 269 -125
rect 273 -123 295 -121
rect 273 -125 284 -123
rect 286 -125 291 -123
rect 293 -125 295 -123
rect 273 -127 295 -125
rect 299 -123 305 -121
rect 299 -125 301 -123
rect 303 -125 305 -123
rect 299 -127 305 -125
rect 309 -123 315 -121
rect 309 -125 311 -123
rect 313 -125 315 -123
rect 309 -127 315 -125
rect 332 -122 338 -120
rect 332 -124 334 -122
rect 336 -124 338 -122
rect 332 -126 338 -124
rect 263 -130 265 -127
rect 273 -130 275 -127
rect 293 -130 295 -127
rect 300 -130 302 -127
rect 191 -149 193 -144
rect 201 -149 203 -144
rect 153 -154 155 -150
rect 164 -154 166 -150
rect 171 -154 173 -150
rect 211 -152 213 -147
rect 221 -154 223 -150
rect 243 -154 245 -150
rect 253 -152 255 -147
rect 263 -149 265 -144
rect 273 -149 275 -144
rect 311 -136 313 -127
rect 332 -135 334 -126
rect 342 -135 344 -119
rect 352 -121 354 -108
rect 395 -93 397 -88
rect 402 -93 404 -88
rect 420 -90 422 -86
rect 430 -90 432 -86
rect 440 -90 442 -86
rect 462 -90 464 -86
rect 472 -90 474 -86
rect 482 -90 484 -86
rect 385 -102 387 -97
rect 352 -123 358 -121
rect 352 -125 354 -123
rect 356 -125 358 -123
rect 352 -127 358 -125
rect 352 -135 354 -127
rect 372 -128 374 -115
rect 385 -118 387 -115
rect 500 -93 502 -88
rect 507 -93 509 -88
rect 530 -90 532 -86
rect 550 -90 552 -86
rect 557 -90 559 -86
rect 517 -102 519 -97
rect 591 -90 593 -86
rect 601 -90 603 -86
rect 611 -90 613 -86
rect 570 -99 572 -95
rect 517 -118 519 -115
rect 378 -120 387 -118
rect 378 -122 380 -120
rect 382 -122 384 -120
rect 395 -121 397 -118
rect 402 -121 404 -118
rect 420 -121 422 -118
rect 430 -121 432 -118
rect 440 -121 442 -118
rect 462 -121 464 -118
rect 472 -121 474 -118
rect 482 -121 484 -118
rect 500 -121 502 -118
rect 507 -121 509 -118
rect 517 -120 526 -118
rect 378 -124 384 -122
rect 372 -130 378 -128
rect 372 -132 374 -130
rect 376 -132 378 -130
rect 372 -134 378 -132
rect 372 -137 374 -134
rect 382 -137 384 -124
rect 392 -123 398 -121
rect 392 -125 394 -123
rect 396 -125 398 -123
rect 392 -127 398 -125
rect 402 -123 424 -121
rect 402 -125 413 -123
rect 415 -125 420 -123
rect 422 -125 424 -123
rect 402 -127 424 -125
rect 428 -123 434 -121
rect 428 -125 430 -123
rect 432 -125 434 -123
rect 428 -127 434 -125
rect 438 -123 444 -121
rect 438 -125 440 -123
rect 442 -125 444 -123
rect 438 -127 444 -125
rect 460 -123 466 -121
rect 460 -125 462 -123
rect 464 -125 466 -123
rect 460 -127 466 -125
rect 470 -123 476 -121
rect 470 -125 472 -123
rect 474 -125 476 -123
rect 470 -127 476 -125
rect 480 -123 502 -121
rect 480 -125 482 -123
rect 484 -125 489 -123
rect 491 -125 502 -123
rect 480 -127 502 -125
rect 506 -123 512 -121
rect 506 -125 508 -123
rect 510 -125 512 -123
rect 506 -127 512 -125
rect 392 -130 394 -127
rect 402 -130 404 -127
rect 422 -130 424 -127
rect 429 -130 431 -127
rect 332 -145 334 -141
rect 342 -145 344 -141
rect 352 -145 354 -141
rect 293 -154 295 -150
rect 300 -154 302 -150
rect 311 -154 313 -150
rect 372 -154 374 -150
rect 382 -152 384 -147
rect 392 -149 394 -144
rect 402 -149 404 -144
rect 440 -136 442 -127
rect 462 -136 464 -127
rect 473 -130 475 -127
rect 480 -130 482 -127
rect 500 -130 502 -127
rect 510 -130 512 -127
rect 520 -122 522 -120
rect 524 -122 526 -120
rect 520 -124 526 -122
rect 520 -137 522 -124
rect 530 -128 532 -115
rect 550 -121 552 -108
rect 557 -113 559 -108
rect 556 -115 562 -113
rect 556 -117 558 -115
rect 560 -117 562 -115
rect 556 -119 562 -117
rect 546 -123 552 -121
rect 546 -125 548 -123
rect 550 -125 552 -123
rect 546 -127 552 -125
rect 526 -130 532 -128
rect 526 -132 528 -130
rect 530 -132 532 -130
rect 526 -134 532 -132
rect 530 -137 532 -134
rect 550 -135 552 -127
rect 560 -135 562 -119
rect 570 -120 572 -111
rect 629 -93 631 -88
rect 636 -93 638 -88
rect 659 -90 661 -86
rect 683 -90 685 -86
rect 693 -90 695 -86
rect 703 -90 705 -86
rect 646 -102 648 -97
rect 646 -118 648 -115
rect 566 -122 572 -120
rect 591 -121 593 -118
rect 601 -121 603 -118
rect 611 -121 613 -118
rect 629 -121 631 -118
rect 636 -121 638 -118
rect 646 -120 655 -118
rect 566 -124 568 -122
rect 570 -124 572 -122
rect 566 -126 572 -124
rect 570 -135 572 -126
rect 589 -123 595 -121
rect 589 -125 591 -123
rect 593 -125 595 -123
rect 589 -127 595 -125
rect 599 -123 605 -121
rect 599 -125 601 -123
rect 603 -125 605 -123
rect 599 -127 605 -125
rect 609 -123 631 -121
rect 609 -125 611 -123
rect 613 -125 618 -123
rect 620 -125 631 -123
rect 609 -127 631 -125
rect 635 -123 641 -121
rect 635 -125 637 -123
rect 639 -125 641 -123
rect 635 -127 641 -125
rect 500 -149 502 -144
rect 510 -149 512 -144
rect 422 -154 424 -150
rect 429 -154 431 -150
rect 440 -154 442 -150
rect 462 -154 464 -150
rect 473 -154 475 -150
rect 480 -154 482 -150
rect 520 -152 522 -147
rect 591 -136 593 -127
rect 602 -130 604 -127
rect 609 -130 611 -127
rect 629 -130 631 -127
rect 639 -130 641 -127
rect 649 -122 651 -120
rect 653 -122 655 -120
rect 649 -124 655 -122
rect 550 -145 552 -141
rect 560 -145 562 -141
rect 570 -145 572 -141
rect 530 -154 532 -150
rect 649 -137 651 -124
rect 659 -128 661 -115
rect 721 -93 723 -88
rect 728 -93 730 -88
rect 751 -90 753 -86
rect 738 -102 740 -97
rect 738 -118 740 -115
rect 683 -121 685 -118
rect 693 -121 695 -118
rect 703 -121 705 -118
rect 721 -121 723 -118
rect 728 -121 730 -118
rect 738 -120 747 -118
rect 681 -123 687 -121
rect 681 -125 683 -123
rect 685 -125 687 -123
rect 681 -127 687 -125
rect 691 -123 697 -121
rect 691 -125 693 -123
rect 695 -125 697 -123
rect 691 -127 697 -125
rect 701 -123 723 -121
rect 701 -125 703 -123
rect 705 -125 710 -123
rect 712 -125 723 -123
rect 701 -127 723 -125
rect 727 -123 733 -121
rect 727 -125 729 -123
rect 731 -125 733 -123
rect 727 -127 733 -125
rect 655 -130 661 -128
rect 655 -132 657 -130
rect 659 -132 661 -130
rect 655 -134 661 -132
rect 659 -137 661 -134
rect 683 -136 685 -127
rect 694 -130 696 -127
rect 701 -130 703 -127
rect 721 -130 723 -127
rect 731 -130 733 -127
rect 741 -122 743 -120
rect 745 -122 747 -120
rect 741 -124 747 -122
rect 629 -149 631 -144
rect 639 -149 641 -144
rect 591 -154 593 -150
rect 602 -154 604 -150
rect 609 -154 611 -150
rect 649 -152 651 -147
rect 741 -137 743 -124
rect 751 -128 753 -115
rect 747 -130 753 -128
rect 747 -132 749 -130
rect 751 -132 753 -130
rect 747 -134 753 -132
rect 751 -137 753 -134
rect 721 -149 723 -144
rect 731 -149 733 -144
rect 659 -154 661 -150
rect 683 -154 685 -150
rect 694 -154 696 -150
rect 701 -154 703 -150
rect 741 -152 743 -147
rect 751 -154 753 -150
rect 438 -231 464 -229
rect 470 -231 550 -229
rect 417 -233 423 -231
rect 417 -235 419 -233
rect 421 -235 423 -233
rect 407 -240 409 -235
rect 417 -237 423 -235
rect 438 -237 440 -231
rect 460 -233 466 -231
rect 460 -235 462 -233
rect 464 -235 466 -233
rect 417 -242 419 -237
rect 427 -239 440 -237
rect 427 -242 429 -239
rect 450 -240 452 -235
rect 460 -237 466 -235
rect 460 -242 462 -237
rect 470 -242 472 -231
rect 546 -233 552 -231
rect 546 -235 548 -233
rect 550 -235 552 -233
rect 493 -240 495 -235
rect 503 -242 505 -238
rect 513 -242 515 -237
rect 536 -240 538 -235
rect 546 -237 552 -235
rect 828 -237 830 178
rect 546 -242 548 -237
rect 556 -239 830 -237
rect 556 -242 558 -239
rect 407 -255 409 -252
rect 417 -255 419 -252
rect 407 -257 413 -255
rect 407 -259 409 -257
rect 411 -259 413 -257
rect 417 -258 421 -255
rect 407 -261 413 -259
rect 407 -269 409 -261
rect 419 -272 421 -258
rect 427 -263 429 -252
rect 450 -255 452 -252
rect 460 -255 462 -252
rect 450 -257 456 -255
rect 450 -259 452 -257
rect 454 -259 456 -257
rect 460 -258 464 -255
rect 450 -261 456 -259
rect 426 -265 432 -263
rect 426 -267 428 -265
rect 430 -267 432 -265
rect 426 -269 432 -267
rect 450 -269 452 -261
rect 426 -272 428 -269
rect 407 -279 409 -275
rect 462 -272 464 -258
rect 470 -263 472 -252
rect 493 -255 495 -252
rect 503 -255 505 -252
rect 493 -257 499 -255
rect 493 -259 495 -257
rect 497 -259 499 -257
rect 503 -258 507 -255
rect 493 -261 499 -259
rect 469 -265 475 -263
rect 469 -267 471 -265
rect 473 -267 475 -265
rect 469 -269 475 -267
rect 493 -269 495 -261
rect 469 -272 471 -269
rect 450 -279 452 -275
rect 505 -272 507 -258
rect 513 -263 515 -252
rect 536 -255 538 -252
rect 546 -255 548 -252
rect 536 -257 542 -255
rect 536 -259 538 -257
rect 540 -259 542 -257
rect 546 -258 550 -255
rect 536 -261 542 -259
rect 512 -265 518 -263
rect 512 -267 514 -265
rect 516 -267 518 -265
rect 512 -269 518 -267
rect 536 -269 538 -261
rect 512 -272 514 -269
rect 493 -279 495 -275
rect 548 -272 550 -258
rect 556 -263 558 -252
rect 555 -265 561 -263
rect 555 -267 557 -265
rect 559 -267 561 -265
rect 555 -269 561 -267
rect 555 -272 557 -269
rect 536 -279 538 -275
rect 419 -293 421 -281
rect 426 -286 428 -281
rect 462 -286 464 -281
rect 469 -286 471 -281
rect 505 -293 507 -281
rect 512 -293 514 -281
rect 548 -286 550 -281
rect 555 -293 557 -281
rect 419 -295 508 -293
rect 512 -295 557 -293
rect 588 -305 596 -301
rect 848 -305 850 202
rect 588 -306 850 -305
rect 588 -308 591 -306
rect 593 -307 850 -306
rect 593 -308 596 -307
rect 588 -311 596 -308
rect 406 -320 408 -316
rect 429 -323 431 -318
rect 436 -323 438 -318
rect 454 -320 456 -316
rect 464 -320 466 -316
rect 474 -320 476 -316
rect 508 -320 510 -316
rect 518 -320 520 -316
rect 528 -320 530 -316
rect 419 -332 421 -327
rect 406 -358 408 -345
rect 419 -348 421 -345
rect 546 -323 548 -318
rect 553 -323 555 -318
rect 576 -320 578 -316
rect 563 -332 565 -327
rect 563 -348 565 -345
rect 412 -350 421 -348
rect 412 -352 414 -350
rect 416 -352 418 -350
rect 429 -351 431 -348
rect 436 -351 438 -348
rect 454 -351 456 -348
rect 464 -351 466 -348
rect 474 -351 476 -348
rect 508 -351 510 -348
rect 518 -351 520 -348
rect 528 -351 530 -348
rect 546 -351 548 -348
rect 553 -351 555 -348
rect 563 -350 572 -348
rect 412 -354 418 -352
rect 406 -360 412 -358
rect 406 -362 408 -360
rect 410 -362 412 -360
rect 406 -364 412 -362
rect 406 -367 408 -364
rect 416 -367 418 -354
rect 426 -353 432 -351
rect 426 -355 428 -353
rect 430 -355 432 -353
rect 426 -357 432 -355
rect 436 -353 458 -351
rect 436 -355 447 -353
rect 449 -355 454 -353
rect 456 -355 458 -353
rect 436 -357 458 -355
rect 462 -353 468 -351
rect 462 -355 464 -353
rect 466 -355 468 -353
rect 462 -357 468 -355
rect 472 -353 478 -351
rect 472 -355 474 -353
rect 476 -355 478 -353
rect 472 -357 478 -355
rect 506 -353 512 -351
rect 506 -355 508 -353
rect 510 -355 512 -353
rect 506 -357 512 -355
rect 516 -353 522 -351
rect 516 -355 518 -353
rect 520 -355 522 -353
rect 516 -357 522 -355
rect 526 -353 548 -351
rect 526 -355 528 -353
rect 530 -355 535 -353
rect 537 -355 548 -353
rect 526 -357 548 -355
rect 552 -353 558 -351
rect 552 -355 554 -353
rect 556 -355 558 -353
rect 552 -357 558 -355
rect 426 -360 428 -357
rect 436 -360 438 -357
rect 456 -360 458 -357
rect 463 -360 465 -357
rect -146 -379 -40 -377
rect 406 -384 408 -380
rect 416 -382 418 -377
rect 426 -379 428 -374
rect 436 -379 438 -374
rect 474 -366 476 -357
rect 508 -366 510 -357
rect 519 -360 521 -357
rect 526 -360 528 -357
rect 546 -360 548 -357
rect 556 -360 558 -357
rect 566 -352 568 -350
rect 570 -352 572 -350
rect 566 -354 572 -352
rect 566 -367 568 -354
rect 576 -358 578 -345
rect 572 -360 578 -358
rect 572 -362 574 -360
rect 576 -362 578 -360
rect 572 -364 578 -362
rect 576 -367 578 -364
rect 546 -379 548 -374
rect 556 -379 558 -374
rect 456 -384 458 -380
rect 463 -384 465 -380
rect 474 -384 476 -380
rect 508 -384 510 -380
rect 519 -384 521 -380
rect 526 -384 528 -380
rect 566 -382 568 -377
rect 576 -384 578 -380
rect -246 -397 -244 -393
rect -223 -400 -221 -395
rect -216 -400 -214 -395
rect -198 -397 -196 -393
rect -188 -397 -186 -393
rect -178 -397 -176 -393
rect -144 -397 -142 -393
rect -134 -397 -132 -393
rect -124 -397 -122 -393
rect -233 -409 -231 -404
rect -246 -435 -244 -422
rect -233 -425 -231 -422
rect -106 -400 -104 -395
rect -99 -400 -97 -395
rect -76 -397 -74 -393
rect -89 -409 -87 -404
rect -89 -425 -87 -422
rect -240 -427 -231 -425
rect -240 -429 -238 -427
rect -236 -429 -234 -427
rect -223 -428 -221 -425
rect -216 -428 -214 -425
rect -198 -428 -196 -425
rect -188 -428 -186 -425
rect -178 -428 -176 -425
rect -144 -428 -142 -425
rect -134 -428 -132 -425
rect -124 -428 -122 -425
rect -106 -428 -104 -425
rect -99 -428 -97 -425
rect -89 -427 -80 -425
rect -240 -431 -234 -429
rect -246 -437 -240 -435
rect -246 -439 -244 -437
rect -242 -439 -240 -437
rect -246 -441 -240 -439
rect -246 -444 -244 -441
rect -236 -444 -234 -431
rect -226 -430 -220 -428
rect -226 -432 -224 -430
rect -222 -432 -220 -430
rect -226 -434 -220 -432
rect -216 -430 -194 -428
rect -216 -432 -205 -430
rect -203 -432 -198 -430
rect -196 -432 -194 -430
rect -216 -434 -194 -432
rect -190 -430 -184 -428
rect -190 -432 -188 -430
rect -186 -432 -184 -430
rect -190 -434 -184 -432
rect -180 -430 -174 -428
rect -180 -432 -178 -430
rect -176 -432 -174 -430
rect -180 -434 -174 -432
rect -146 -430 -140 -428
rect -146 -432 -144 -430
rect -142 -432 -140 -430
rect -146 -434 -140 -432
rect -136 -430 -130 -428
rect -136 -432 -134 -430
rect -132 -432 -130 -430
rect -136 -434 -130 -432
rect -126 -430 -104 -428
rect -126 -432 -124 -430
rect -122 -432 -117 -430
rect -115 -432 -104 -430
rect -126 -434 -104 -432
rect -100 -430 -94 -428
rect -100 -432 -98 -430
rect -96 -432 -94 -430
rect -100 -434 -94 -432
rect -226 -437 -224 -434
rect -216 -437 -214 -434
rect -196 -437 -194 -434
rect -189 -437 -187 -434
rect -246 -461 -244 -457
rect -236 -458 -234 -454
rect -226 -456 -224 -451
rect -216 -456 -214 -451
rect -178 -443 -176 -434
rect -144 -443 -142 -434
rect -133 -437 -131 -434
rect -126 -437 -124 -434
rect -106 -437 -104 -434
rect -96 -437 -94 -434
rect -86 -429 -84 -427
rect -82 -429 -80 -427
rect -86 -431 -80 -429
rect -86 -444 -84 -431
rect -76 -435 -74 -422
rect -80 -437 -74 -435
rect -80 -439 -78 -437
rect -76 -439 -74 -437
rect -80 -441 -74 -439
rect -76 -444 -74 -441
rect -106 -456 -104 -451
rect -96 -456 -94 -451
rect -196 -461 -194 -457
rect -189 -461 -187 -457
rect -178 -461 -176 -457
rect -144 -461 -142 -457
rect -133 -461 -131 -457
rect -126 -461 -124 -457
rect -86 -459 -84 -454
rect -76 -461 -74 -457
rect 26 -475 28 -471
rect 36 -475 38 -471
rect 46 -475 48 -471
rect 64 -478 66 -473
rect 71 -478 73 -473
rect 94 -475 96 -471
rect 114 -475 116 -471
rect 121 -475 123 -471
rect 81 -487 83 -482
rect 155 -475 157 -471
rect 165 -475 167 -471
rect 175 -475 177 -471
rect 134 -484 136 -480
rect 81 -503 83 -500
rect 26 -506 28 -503
rect 36 -506 38 -503
rect 46 -506 48 -503
rect 64 -506 66 -503
rect 71 -506 73 -503
rect 81 -505 90 -503
rect 24 -508 30 -506
rect 24 -510 26 -508
rect 28 -510 30 -508
rect 24 -512 30 -510
rect 34 -508 40 -506
rect 34 -510 36 -508
rect 38 -510 40 -508
rect 34 -512 40 -510
rect 44 -508 66 -506
rect 44 -510 46 -508
rect 48 -510 53 -508
rect 55 -510 66 -508
rect 44 -512 66 -510
rect 70 -508 76 -506
rect 70 -510 72 -508
rect 74 -510 76 -508
rect 70 -512 76 -510
rect 26 -521 28 -512
rect 37 -515 39 -512
rect 44 -515 46 -512
rect 64 -515 66 -512
rect 74 -515 76 -512
rect 84 -507 86 -505
rect 88 -507 90 -505
rect 84 -509 90 -507
rect 84 -522 86 -509
rect 94 -513 96 -500
rect 114 -506 116 -493
rect 121 -498 123 -493
rect 120 -500 126 -498
rect 120 -502 122 -500
rect 124 -502 126 -500
rect 120 -504 126 -502
rect 110 -508 116 -506
rect 110 -510 112 -508
rect 114 -510 116 -508
rect 110 -512 116 -510
rect 90 -515 96 -513
rect 90 -517 92 -515
rect 94 -517 96 -515
rect 90 -519 96 -517
rect 94 -522 96 -519
rect 114 -520 116 -512
rect 124 -520 126 -504
rect 134 -505 136 -496
rect 193 -478 195 -473
rect 200 -478 202 -473
rect 223 -475 225 -471
rect 245 -475 247 -471
rect 210 -487 212 -482
rect 268 -478 270 -473
rect 275 -478 277 -473
rect 293 -475 295 -471
rect 303 -475 305 -471
rect 313 -475 315 -471
rect 258 -487 260 -482
rect 210 -503 212 -500
rect 130 -507 136 -505
rect 155 -506 157 -503
rect 165 -506 167 -503
rect 175 -506 177 -503
rect 193 -506 195 -503
rect 200 -506 202 -503
rect 210 -505 219 -503
rect 130 -509 132 -507
rect 134 -509 136 -507
rect 130 -511 136 -509
rect 134 -520 136 -511
rect 153 -508 159 -506
rect 153 -510 155 -508
rect 157 -510 159 -508
rect 153 -512 159 -510
rect 163 -508 169 -506
rect 163 -510 165 -508
rect 167 -510 169 -508
rect 163 -512 169 -510
rect 173 -508 195 -506
rect 173 -510 175 -508
rect 177 -510 182 -508
rect 184 -510 195 -508
rect 173 -512 195 -510
rect 199 -508 205 -506
rect 199 -510 201 -508
rect 203 -510 205 -508
rect 199 -512 205 -510
rect 64 -534 66 -529
rect 74 -534 76 -529
rect 26 -539 28 -535
rect 37 -539 39 -535
rect 44 -539 46 -535
rect 84 -537 86 -532
rect 155 -521 157 -512
rect 166 -515 168 -512
rect 173 -515 175 -512
rect 193 -515 195 -512
rect 203 -515 205 -512
rect 213 -507 215 -505
rect 217 -507 219 -505
rect 213 -509 219 -507
rect 114 -530 116 -526
rect 124 -530 126 -526
rect 134 -530 136 -526
rect 94 -539 96 -535
rect 213 -522 215 -509
rect 223 -513 225 -500
rect 219 -515 225 -513
rect 219 -517 221 -515
rect 223 -517 225 -515
rect 219 -519 225 -517
rect 223 -522 225 -519
rect 245 -513 247 -500
rect 258 -503 260 -500
rect 347 -475 349 -471
rect 354 -475 356 -471
rect 374 -475 376 -471
rect 334 -484 336 -480
rect 251 -505 260 -503
rect 251 -507 253 -505
rect 255 -507 257 -505
rect 268 -506 270 -503
rect 275 -506 277 -503
rect 293 -506 295 -503
rect 303 -506 305 -503
rect 313 -506 315 -503
rect 334 -505 336 -496
rect 347 -498 349 -493
rect 344 -500 350 -498
rect 344 -502 346 -500
rect 348 -502 350 -500
rect 344 -504 350 -502
rect 251 -509 257 -507
rect 245 -515 251 -513
rect 245 -517 247 -515
rect 249 -517 251 -515
rect 245 -519 251 -517
rect 245 -522 247 -519
rect 255 -522 257 -509
rect 265 -508 271 -506
rect 265 -510 267 -508
rect 269 -510 271 -508
rect 265 -512 271 -510
rect 275 -508 297 -506
rect 275 -510 286 -508
rect 288 -510 293 -508
rect 295 -510 297 -508
rect 275 -512 297 -510
rect 301 -508 307 -506
rect 301 -510 303 -508
rect 305 -510 307 -508
rect 301 -512 307 -510
rect 311 -508 317 -506
rect 311 -510 313 -508
rect 315 -510 317 -508
rect 311 -512 317 -510
rect 334 -507 340 -505
rect 334 -509 336 -507
rect 338 -509 340 -507
rect 334 -511 340 -509
rect 265 -515 267 -512
rect 275 -515 277 -512
rect 295 -515 297 -512
rect 302 -515 304 -512
rect 193 -534 195 -529
rect 203 -534 205 -529
rect 155 -539 157 -535
rect 166 -539 168 -535
rect 173 -539 175 -535
rect 213 -537 215 -532
rect 223 -539 225 -535
rect 245 -539 247 -535
rect 255 -537 257 -532
rect 265 -534 267 -529
rect 275 -534 277 -529
rect 313 -521 315 -512
rect 334 -520 336 -511
rect 344 -520 346 -504
rect 354 -506 356 -493
rect 397 -478 399 -473
rect 404 -478 406 -473
rect 422 -475 424 -471
rect 432 -475 434 -471
rect 442 -475 444 -471
rect 464 -475 466 -471
rect 474 -475 476 -471
rect 484 -475 486 -471
rect 387 -487 389 -482
rect 354 -508 360 -506
rect 354 -510 356 -508
rect 358 -510 360 -508
rect 354 -512 360 -510
rect 354 -520 356 -512
rect 374 -513 376 -500
rect 387 -503 389 -500
rect 502 -478 504 -473
rect 509 -478 511 -473
rect 532 -475 534 -471
rect 552 -475 554 -471
rect 559 -475 561 -471
rect 519 -487 521 -482
rect 593 -475 595 -471
rect 603 -475 605 -471
rect 613 -475 615 -471
rect 572 -484 574 -480
rect 519 -503 521 -500
rect 380 -505 389 -503
rect 380 -507 382 -505
rect 384 -507 386 -505
rect 397 -506 399 -503
rect 404 -506 406 -503
rect 422 -506 424 -503
rect 432 -506 434 -503
rect 442 -506 444 -503
rect 464 -506 466 -503
rect 474 -506 476 -503
rect 484 -506 486 -503
rect 502 -506 504 -503
rect 509 -506 511 -503
rect 519 -505 528 -503
rect 380 -509 386 -507
rect 374 -515 380 -513
rect 374 -517 376 -515
rect 378 -517 380 -515
rect 374 -519 380 -517
rect 374 -522 376 -519
rect 384 -522 386 -509
rect 394 -508 400 -506
rect 394 -510 396 -508
rect 398 -510 400 -508
rect 394 -512 400 -510
rect 404 -508 426 -506
rect 404 -510 415 -508
rect 417 -510 422 -508
rect 424 -510 426 -508
rect 404 -512 426 -510
rect 430 -508 436 -506
rect 430 -510 432 -508
rect 434 -510 436 -508
rect 430 -512 436 -510
rect 440 -508 446 -506
rect 440 -510 442 -508
rect 444 -510 446 -508
rect 440 -512 446 -510
rect 462 -508 468 -506
rect 462 -510 464 -508
rect 466 -510 468 -508
rect 462 -512 468 -510
rect 472 -508 478 -506
rect 472 -510 474 -508
rect 476 -510 478 -508
rect 472 -512 478 -510
rect 482 -508 504 -506
rect 482 -510 484 -508
rect 486 -510 491 -508
rect 493 -510 504 -508
rect 482 -512 504 -510
rect 508 -508 514 -506
rect 508 -510 510 -508
rect 512 -510 514 -508
rect 508 -512 514 -510
rect 394 -515 396 -512
rect 404 -515 406 -512
rect 424 -515 426 -512
rect 431 -515 433 -512
rect 334 -530 336 -526
rect 344 -530 346 -526
rect 354 -530 356 -526
rect 295 -539 297 -535
rect 302 -539 304 -535
rect 313 -539 315 -535
rect 374 -539 376 -535
rect 384 -537 386 -532
rect 394 -534 396 -529
rect 404 -534 406 -529
rect 442 -521 444 -512
rect 464 -521 466 -512
rect 475 -515 477 -512
rect 482 -515 484 -512
rect 502 -515 504 -512
rect 512 -515 514 -512
rect 522 -507 524 -505
rect 526 -507 528 -505
rect 522 -509 528 -507
rect 522 -522 524 -509
rect 532 -513 534 -500
rect 552 -506 554 -493
rect 559 -498 561 -493
rect 558 -500 564 -498
rect 558 -502 560 -500
rect 562 -502 564 -500
rect 558 -504 564 -502
rect 548 -508 554 -506
rect 548 -510 550 -508
rect 552 -510 554 -508
rect 548 -512 554 -510
rect 528 -515 534 -513
rect 528 -517 530 -515
rect 532 -517 534 -515
rect 528 -519 534 -517
rect 532 -522 534 -519
rect 552 -520 554 -512
rect 562 -520 564 -504
rect 572 -505 574 -496
rect 631 -478 633 -473
rect 638 -478 640 -473
rect 661 -475 663 -471
rect 685 -475 687 -471
rect 695 -475 697 -471
rect 705 -475 707 -471
rect 648 -487 650 -482
rect 648 -503 650 -500
rect 568 -507 574 -505
rect 593 -506 595 -503
rect 603 -506 605 -503
rect 613 -506 615 -503
rect 631 -506 633 -503
rect 638 -506 640 -503
rect 648 -505 657 -503
rect 568 -509 570 -507
rect 572 -509 574 -507
rect 568 -511 574 -509
rect 572 -520 574 -511
rect 591 -508 597 -506
rect 591 -510 593 -508
rect 595 -510 597 -508
rect 591 -512 597 -510
rect 601 -508 607 -506
rect 601 -510 603 -508
rect 605 -510 607 -508
rect 601 -512 607 -510
rect 611 -508 633 -506
rect 611 -510 613 -508
rect 615 -510 620 -508
rect 622 -510 633 -508
rect 611 -512 633 -510
rect 637 -508 643 -506
rect 637 -510 639 -508
rect 641 -510 643 -508
rect 637 -512 643 -510
rect 502 -534 504 -529
rect 512 -534 514 -529
rect 424 -539 426 -535
rect 431 -539 433 -535
rect 442 -539 444 -535
rect 464 -539 466 -535
rect 475 -539 477 -535
rect 482 -539 484 -535
rect 522 -537 524 -532
rect 593 -521 595 -512
rect 604 -515 606 -512
rect 611 -515 613 -512
rect 631 -515 633 -512
rect 641 -515 643 -512
rect 651 -507 653 -505
rect 655 -507 657 -505
rect 651 -509 657 -507
rect 552 -530 554 -526
rect 562 -530 564 -526
rect 572 -530 574 -526
rect 532 -539 534 -535
rect 651 -522 653 -509
rect 661 -513 663 -500
rect 723 -478 725 -473
rect 730 -478 732 -473
rect 753 -475 755 -471
rect 740 -487 742 -482
rect 740 -503 742 -500
rect 685 -506 687 -503
rect 695 -506 697 -503
rect 705 -506 707 -503
rect 723 -506 725 -503
rect 730 -506 732 -503
rect 740 -505 749 -503
rect 683 -508 689 -506
rect 683 -510 685 -508
rect 687 -510 689 -508
rect 683 -512 689 -510
rect 693 -508 699 -506
rect 693 -510 695 -508
rect 697 -510 699 -508
rect 693 -512 699 -510
rect 703 -508 725 -506
rect 703 -510 705 -508
rect 707 -510 712 -508
rect 714 -510 725 -508
rect 703 -512 725 -510
rect 729 -508 735 -506
rect 729 -510 731 -508
rect 733 -510 735 -508
rect 729 -512 735 -510
rect 657 -515 663 -513
rect 657 -517 659 -515
rect 661 -517 663 -515
rect 657 -519 663 -517
rect 661 -522 663 -519
rect 685 -521 687 -512
rect 696 -515 698 -512
rect 703 -515 705 -512
rect 723 -515 725 -512
rect 733 -515 735 -512
rect 743 -507 745 -505
rect 747 -507 749 -505
rect 743 -509 749 -507
rect 631 -534 633 -529
rect 641 -534 643 -529
rect 593 -539 595 -535
rect 604 -539 606 -535
rect 611 -539 613 -535
rect 651 -537 653 -532
rect 743 -522 745 -509
rect 753 -513 755 -500
rect 749 -515 755 -513
rect 749 -517 751 -515
rect 753 -517 755 -515
rect 749 -519 755 -517
rect 753 -522 755 -519
rect 723 -534 725 -529
rect 733 -534 735 -529
rect 661 -539 663 -535
rect 685 -539 687 -535
rect 696 -539 698 -535
rect 703 -539 705 -535
rect 743 -537 745 -532
rect 753 -539 755 -535
rect -241 -609 -239 -605
rect -231 -609 -229 -605
rect -221 -609 -219 -605
rect -203 -612 -201 -607
rect -196 -612 -194 -607
rect -173 -609 -171 -605
rect -153 -609 -151 -605
rect -146 -609 -144 -605
rect -186 -621 -184 -616
rect -112 -609 -110 -605
rect -102 -609 -100 -605
rect -92 -609 -90 -605
rect -133 -618 -131 -614
rect -186 -637 -184 -634
rect -241 -640 -239 -637
rect -231 -640 -229 -637
rect -221 -640 -219 -637
rect -203 -640 -201 -637
rect -196 -640 -194 -637
rect -186 -639 -177 -637
rect -243 -642 -237 -640
rect -243 -644 -241 -642
rect -239 -644 -237 -642
rect -243 -646 -237 -644
rect -233 -642 -227 -640
rect -233 -644 -231 -642
rect -229 -644 -227 -642
rect -233 -646 -227 -644
rect -223 -642 -201 -640
rect -223 -644 -221 -642
rect -219 -644 -214 -642
rect -212 -644 -201 -642
rect -223 -646 -201 -644
rect -197 -642 -191 -640
rect -197 -644 -195 -642
rect -193 -644 -191 -642
rect -197 -646 -191 -644
rect -241 -655 -239 -646
rect -230 -649 -228 -646
rect -223 -649 -221 -646
rect -203 -649 -201 -646
rect -193 -649 -191 -646
rect -183 -641 -181 -639
rect -179 -641 -177 -639
rect -183 -643 -177 -641
rect -183 -656 -181 -643
rect -173 -647 -171 -634
rect -153 -640 -151 -627
rect -146 -632 -144 -627
rect -147 -634 -141 -632
rect -147 -636 -145 -634
rect -143 -636 -141 -634
rect -147 -638 -141 -636
rect -157 -642 -151 -640
rect -157 -644 -155 -642
rect -153 -644 -151 -642
rect -157 -646 -151 -644
rect -177 -649 -171 -647
rect -177 -651 -175 -649
rect -173 -651 -171 -649
rect -177 -653 -171 -651
rect -173 -656 -171 -653
rect -153 -654 -151 -646
rect -143 -654 -141 -638
rect -133 -639 -131 -630
rect -74 -612 -72 -607
rect -67 -612 -65 -607
rect -44 -609 -42 -605
rect -22 -609 -20 -605
rect -57 -621 -55 -616
rect 1 -612 3 -607
rect 8 -612 10 -607
rect 26 -609 28 -605
rect 36 -609 38 -605
rect 46 -609 48 -605
rect -9 -621 -7 -616
rect -57 -637 -55 -634
rect -137 -641 -131 -639
rect -112 -640 -110 -637
rect -102 -640 -100 -637
rect -92 -640 -90 -637
rect -74 -640 -72 -637
rect -67 -640 -65 -637
rect -57 -639 -48 -637
rect -137 -643 -135 -641
rect -133 -643 -131 -641
rect -137 -645 -131 -643
rect -133 -654 -131 -645
rect -114 -642 -108 -640
rect -114 -644 -112 -642
rect -110 -644 -108 -642
rect -114 -646 -108 -644
rect -104 -642 -98 -640
rect -104 -644 -102 -642
rect -100 -644 -98 -642
rect -104 -646 -98 -644
rect -94 -642 -72 -640
rect -94 -644 -92 -642
rect -90 -644 -85 -642
rect -83 -644 -72 -642
rect -94 -646 -72 -644
rect -68 -642 -62 -640
rect -68 -644 -66 -642
rect -64 -644 -62 -642
rect -68 -646 -62 -644
rect -203 -668 -201 -663
rect -193 -668 -191 -663
rect -241 -673 -239 -669
rect -230 -673 -228 -669
rect -223 -673 -221 -669
rect -183 -671 -181 -666
rect -112 -655 -110 -646
rect -101 -649 -99 -646
rect -94 -649 -92 -646
rect -74 -649 -72 -646
rect -64 -649 -62 -646
rect -54 -641 -52 -639
rect -50 -641 -48 -639
rect -54 -643 -48 -641
rect -153 -664 -151 -660
rect -143 -664 -141 -660
rect -133 -664 -131 -660
rect -173 -673 -171 -669
rect -54 -656 -52 -643
rect -44 -647 -42 -634
rect -48 -649 -42 -647
rect -48 -651 -46 -649
rect -44 -651 -42 -649
rect -48 -653 -42 -651
rect -44 -656 -42 -653
rect -22 -647 -20 -634
rect -9 -637 -7 -634
rect 80 -609 82 -605
rect 87 -609 89 -605
rect 107 -609 109 -605
rect 67 -618 69 -614
rect -16 -639 -7 -637
rect -16 -641 -14 -639
rect -12 -641 -10 -639
rect 1 -640 3 -637
rect 8 -640 10 -637
rect 26 -640 28 -637
rect 36 -640 38 -637
rect 46 -640 48 -637
rect 67 -639 69 -630
rect 80 -632 82 -627
rect 77 -634 83 -632
rect 77 -636 79 -634
rect 81 -636 83 -634
rect 77 -638 83 -636
rect -16 -643 -10 -641
rect -22 -649 -16 -647
rect -22 -651 -20 -649
rect -18 -651 -16 -649
rect -22 -653 -16 -651
rect -22 -656 -20 -653
rect -12 -656 -10 -643
rect -2 -642 4 -640
rect -2 -644 0 -642
rect 2 -644 4 -642
rect -2 -646 4 -644
rect 8 -642 30 -640
rect 8 -644 19 -642
rect 21 -644 26 -642
rect 28 -644 30 -642
rect 8 -646 30 -644
rect 34 -642 40 -640
rect 34 -644 36 -642
rect 38 -644 40 -642
rect 34 -646 40 -644
rect 44 -642 50 -640
rect 44 -644 46 -642
rect 48 -644 50 -642
rect 44 -646 50 -644
rect 67 -641 73 -639
rect 67 -643 69 -641
rect 71 -643 73 -641
rect 67 -645 73 -643
rect -2 -649 0 -646
rect 8 -649 10 -646
rect 28 -649 30 -646
rect 35 -649 37 -646
rect -74 -668 -72 -663
rect -64 -668 -62 -663
rect -112 -673 -110 -669
rect -101 -673 -99 -669
rect -94 -673 -92 -669
rect -54 -671 -52 -666
rect -44 -673 -42 -669
rect -22 -673 -20 -669
rect -12 -671 -10 -666
rect -2 -668 0 -663
rect 8 -668 10 -663
rect 46 -655 48 -646
rect 67 -654 69 -645
rect 77 -654 79 -638
rect 87 -640 89 -627
rect 130 -612 132 -607
rect 137 -612 139 -607
rect 155 -609 157 -605
rect 165 -609 167 -605
rect 175 -609 177 -605
rect 197 -609 199 -605
rect 207 -609 209 -605
rect 217 -609 219 -605
rect 120 -621 122 -616
rect 87 -642 93 -640
rect 87 -644 89 -642
rect 91 -644 93 -642
rect 87 -646 93 -644
rect 87 -654 89 -646
rect 107 -647 109 -634
rect 120 -637 122 -634
rect 235 -612 237 -607
rect 242 -612 244 -607
rect 265 -609 267 -605
rect 285 -609 287 -605
rect 292 -609 294 -605
rect 252 -621 254 -616
rect 326 -609 328 -605
rect 336 -609 338 -605
rect 346 -609 348 -605
rect 305 -618 307 -614
rect 252 -637 254 -634
rect 113 -639 122 -637
rect 113 -641 115 -639
rect 117 -641 119 -639
rect 130 -640 132 -637
rect 137 -640 139 -637
rect 155 -640 157 -637
rect 165 -640 167 -637
rect 175 -640 177 -637
rect 197 -640 199 -637
rect 207 -640 209 -637
rect 217 -640 219 -637
rect 235 -640 237 -637
rect 242 -640 244 -637
rect 252 -639 261 -637
rect 113 -643 119 -641
rect 107 -649 113 -647
rect 107 -651 109 -649
rect 111 -651 113 -649
rect 107 -653 113 -651
rect 107 -656 109 -653
rect 117 -656 119 -643
rect 127 -642 133 -640
rect 127 -644 129 -642
rect 131 -644 133 -642
rect 127 -646 133 -644
rect 137 -642 159 -640
rect 137 -644 148 -642
rect 150 -644 155 -642
rect 157 -644 159 -642
rect 137 -646 159 -644
rect 163 -642 169 -640
rect 163 -644 165 -642
rect 167 -644 169 -642
rect 163 -646 169 -644
rect 173 -642 179 -640
rect 173 -644 175 -642
rect 177 -644 179 -642
rect 173 -646 179 -644
rect 195 -642 201 -640
rect 195 -644 197 -642
rect 199 -644 201 -642
rect 195 -646 201 -644
rect 205 -642 211 -640
rect 205 -644 207 -642
rect 209 -644 211 -642
rect 205 -646 211 -644
rect 215 -642 237 -640
rect 215 -644 217 -642
rect 219 -644 224 -642
rect 226 -644 237 -642
rect 215 -646 237 -644
rect 241 -642 247 -640
rect 241 -644 243 -642
rect 245 -644 247 -642
rect 241 -646 247 -644
rect 127 -649 129 -646
rect 137 -649 139 -646
rect 157 -649 159 -646
rect 164 -649 166 -646
rect 67 -664 69 -660
rect 77 -664 79 -660
rect 87 -664 89 -660
rect 28 -673 30 -669
rect 35 -673 37 -669
rect 46 -673 48 -669
rect 107 -673 109 -669
rect 117 -671 119 -666
rect 127 -668 129 -663
rect 137 -668 139 -663
rect 175 -655 177 -646
rect 197 -655 199 -646
rect 208 -649 210 -646
rect 215 -649 217 -646
rect 235 -649 237 -646
rect 245 -649 247 -646
rect 255 -641 257 -639
rect 259 -641 261 -639
rect 255 -643 261 -641
rect 255 -656 257 -643
rect 265 -647 267 -634
rect 285 -640 287 -627
rect 292 -632 294 -627
rect 291 -634 297 -632
rect 291 -636 293 -634
rect 295 -636 297 -634
rect 291 -638 297 -636
rect 281 -642 287 -640
rect 281 -644 283 -642
rect 285 -644 287 -642
rect 281 -646 287 -644
rect 261 -649 267 -647
rect 261 -651 263 -649
rect 265 -651 267 -649
rect 261 -653 267 -651
rect 265 -656 267 -653
rect 285 -654 287 -646
rect 295 -654 297 -638
rect 305 -639 307 -630
rect 364 -612 366 -607
rect 371 -612 373 -607
rect 394 -609 396 -605
rect 418 -609 420 -605
rect 428 -609 430 -605
rect 438 -609 440 -605
rect 381 -621 383 -616
rect 381 -637 383 -634
rect 301 -641 307 -639
rect 326 -640 328 -637
rect 336 -640 338 -637
rect 346 -640 348 -637
rect 364 -640 366 -637
rect 371 -640 373 -637
rect 381 -639 390 -637
rect 301 -643 303 -641
rect 305 -643 307 -641
rect 301 -645 307 -643
rect 305 -654 307 -645
rect 324 -642 330 -640
rect 324 -644 326 -642
rect 328 -644 330 -642
rect 324 -646 330 -644
rect 334 -642 340 -640
rect 334 -644 336 -642
rect 338 -644 340 -642
rect 334 -646 340 -644
rect 344 -642 366 -640
rect 344 -644 346 -642
rect 348 -644 353 -642
rect 355 -644 366 -642
rect 344 -646 366 -644
rect 370 -642 376 -640
rect 370 -644 372 -642
rect 374 -644 376 -642
rect 370 -646 376 -644
rect 235 -668 237 -663
rect 245 -668 247 -663
rect 157 -673 159 -669
rect 164 -673 166 -669
rect 175 -673 177 -669
rect 197 -673 199 -669
rect 208 -673 210 -669
rect 215 -673 217 -669
rect 255 -671 257 -666
rect 326 -655 328 -646
rect 337 -649 339 -646
rect 344 -649 346 -646
rect 364 -649 366 -646
rect 374 -649 376 -646
rect 384 -641 386 -639
rect 388 -641 390 -639
rect 384 -643 390 -641
rect 285 -664 287 -660
rect 295 -664 297 -660
rect 305 -664 307 -660
rect 265 -673 267 -669
rect 384 -656 386 -643
rect 394 -647 396 -634
rect 456 -612 458 -607
rect 463 -612 465 -607
rect 486 -609 488 -605
rect 473 -621 475 -616
rect 473 -637 475 -634
rect 418 -640 420 -637
rect 428 -640 430 -637
rect 438 -640 440 -637
rect 456 -640 458 -637
rect 463 -640 465 -637
rect 473 -639 482 -637
rect 416 -642 422 -640
rect 416 -644 418 -642
rect 420 -644 422 -642
rect 416 -646 422 -644
rect 426 -642 432 -640
rect 426 -644 428 -642
rect 430 -644 432 -642
rect 426 -646 432 -644
rect 436 -642 458 -640
rect 436 -644 438 -642
rect 440 -644 445 -642
rect 447 -644 458 -642
rect 436 -646 458 -644
rect 462 -642 468 -640
rect 462 -644 464 -642
rect 466 -644 468 -642
rect 462 -646 468 -644
rect 390 -649 396 -647
rect 390 -651 392 -649
rect 394 -651 396 -649
rect 390 -653 396 -651
rect 394 -656 396 -653
rect 418 -655 420 -646
rect 429 -649 431 -646
rect 436 -649 438 -646
rect 456 -649 458 -646
rect 466 -649 468 -646
rect 476 -641 478 -639
rect 480 -641 482 -639
rect 476 -643 482 -641
rect 364 -668 366 -663
rect 374 -668 376 -663
rect 326 -673 328 -669
rect 337 -673 339 -669
rect 344 -673 346 -669
rect 384 -671 386 -666
rect 476 -656 478 -643
rect 486 -647 488 -634
rect 482 -649 488 -647
rect 482 -651 484 -649
rect 486 -651 488 -649
rect 482 -653 488 -651
rect 486 -656 488 -653
rect 456 -668 458 -663
rect 466 -668 468 -663
rect 394 -673 396 -669
rect 418 -673 420 -669
rect 429 -673 431 -669
rect 436 -673 438 -669
rect 476 -671 478 -666
rect 486 -673 488 -669
<< ndif >>
rect -253 -96 -246 -94
rect -253 -98 -251 -96
rect -249 -98 -246 -96
rect -253 -100 -246 -98
rect -244 -97 -236 -94
rect -210 -96 -203 -94
rect -244 -100 -234 -97
rect -242 -106 -234 -100
rect -232 -106 -227 -97
rect -225 -99 -218 -97
rect -225 -101 -222 -99
rect -220 -101 -218 -99
rect -210 -98 -208 -96
rect -206 -98 -203 -96
rect -210 -100 -203 -98
rect -201 -97 -193 -94
rect -167 -96 -160 -94
rect -201 -100 -191 -97
rect -225 -103 -218 -101
rect -225 -106 -220 -103
rect -199 -106 -191 -100
rect -189 -106 -184 -97
rect -182 -99 -175 -97
rect -182 -101 -179 -99
rect -177 -101 -175 -99
rect -167 -98 -165 -96
rect -163 -98 -160 -96
rect -167 -100 -160 -98
rect -158 -97 -150 -94
rect -124 -96 -117 -94
rect -158 -100 -148 -97
rect -182 -103 -175 -101
rect -182 -106 -177 -103
rect -156 -106 -148 -100
rect -146 -106 -141 -97
rect -139 -99 -132 -97
rect -139 -101 -136 -99
rect -134 -101 -132 -99
rect -124 -98 -122 -96
rect -120 -98 -117 -96
rect -124 -100 -117 -98
rect -115 -97 -107 -94
rect -115 -100 -105 -97
rect -139 -103 -132 -101
rect -139 -106 -134 -103
rect -113 -106 -105 -100
rect -103 -106 -98 -97
rect -96 -99 -89 -97
rect -96 -101 -93 -99
rect -91 -101 -89 -99
rect -96 -103 -89 -101
rect -96 -106 -91 -103
rect -242 -108 -236 -106
rect -242 -110 -240 -108
rect -238 -110 -236 -108
rect -242 -112 -236 -110
rect -199 -108 -193 -106
rect -199 -110 -197 -108
rect -195 -110 -193 -108
rect -199 -112 -193 -110
rect -156 -108 -150 -106
rect -156 -110 -154 -108
rect -152 -110 -150 -108
rect -156 -112 -150 -110
rect -113 -108 -107 -106
rect -113 -110 -111 -108
rect -109 -110 -107 -108
rect -113 -112 -107 -110
rect -232 -192 -227 -185
rect -254 -194 -247 -192
rect -254 -196 -252 -194
rect -250 -196 -247 -194
rect -254 -198 -247 -196
rect -252 -205 -247 -198
rect -245 -198 -237 -192
rect -245 -200 -242 -198
rect -240 -200 -237 -198
rect -245 -202 -237 -200
rect -235 -195 -227 -192
rect -235 -197 -232 -195
rect -230 -197 -227 -195
rect -235 -199 -227 -197
rect -225 -187 -217 -185
rect -225 -189 -222 -187
rect -220 -189 -217 -187
rect -225 -199 -217 -189
rect -215 -187 -208 -185
rect -215 -189 -212 -187
rect -210 -189 -208 -187
rect -215 -194 -208 -189
rect -202 -192 -197 -185
rect -215 -196 -212 -194
rect -210 -196 -208 -194
rect -215 -199 -208 -196
rect -204 -194 -197 -192
rect -204 -196 -202 -194
rect -200 -196 -197 -194
rect -204 -198 -197 -196
rect -235 -202 -230 -199
rect -245 -205 -240 -202
rect -202 -205 -197 -198
rect -195 -205 -190 -185
rect -188 -191 -181 -185
rect -141 -191 -134 -185
rect -188 -201 -179 -191
rect -188 -203 -185 -201
rect -183 -203 -179 -201
rect -188 -205 -179 -203
rect -177 -194 -170 -191
rect -177 -196 -174 -194
rect -172 -196 -170 -194
rect -177 -198 -170 -196
rect -152 -194 -145 -191
rect -152 -196 -150 -194
rect -148 -196 -145 -194
rect -152 -198 -145 -196
rect -177 -205 -172 -198
rect -150 -205 -145 -198
rect -143 -201 -134 -191
rect -143 -203 -139 -201
rect -137 -203 -134 -201
rect -143 -205 -134 -203
rect -132 -205 -127 -185
rect -125 -192 -120 -185
rect -114 -187 -107 -185
rect -114 -189 -112 -187
rect -110 -189 -107 -187
rect -125 -194 -118 -192
rect -125 -196 -122 -194
rect -120 -196 -118 -194
rect -125 -198 -118 -196
rect -114 -194 -107 -189
rect -114 -196 -112 -194
rect -110 -196 -107 -194
rect -125 -205 -120 -198
rect -114 -199 -107 -196
rect -105 -187 -97 -185
rect -105 -189 -102 -187
rect -100 -189 -97 -187
rect -105 -199 -97 -189
rect -95 -192 -90 -185
rect -95 -195 -87 -192
rect -95 -197 -92 -195
rect -90 -197 -87 -195
rect -95 -199 -87 -197
rect -92 -202 -87 -199
rect -85 -198 -77 -192
rect -85 -200 -82 -198
rect -80 -200 -77 -198
rect -85 -202 -77 -200
rect -82 -205 -77 -202
rect -75 -194 -68 -192
rect -75 -196 -72 -194
rect -70 -196 -68 -194
rect -75 -198 -68 -196
rect -75 -205 -70 -198
rect -252 -348 -245 -346
rect -252 -350 -250 -348
rect -248 -350 -245 -348
rect -252 -352 -245 -350
rect -243 -349 -235 -346
rect -209 -348 -202 -346
rect -243 -352 -233 -349
rect -241 -358 -233 -352
rect -231 -358 -226 -349
rect -224 -351 -217 -349
rect -224 -353 -221 -351
rect -219 -353 -217 -351
rect -209 -350 -207 -348
rect -205 -350 -202 -348
rect -209 -352 -202 -350
rect -200 -349 -192 -346
rect -166 -348 -159 -346
rect -200 -352 -190 -349
rect -224 -355 -217 -353
rect -224 -358 -219 -355
rect -198 -358 -190 -352
rect -188 -358 -183 -349
rect -181 -351 -174 -349
rect -181 -353 -178 -351
rect -176 -353 -174 -351
rect -166 -350 -164 -348
rect -162 -350 -159 -348
rect -166 -352 -159 -350
rect -157 -349 -149 -346
rect -123 -348 -116 -346
rect -157 -352 -147 -349
rect -181 -355 -174 -353
rect -181 -358 -176 -355
rect -155 -358 -147 -352
rect -145 -358 -140 -349
rect -138 -351 -131 -349
rect -138 -353 -135 -351
rect -133 -353 -131 -351
rect -123 -350 -121 -348
rect -119 -350 -116 -348
rect -123 -352 -116 -350
rect -114 -349 -106 -346
rect -114 -352 -104 -349
rect -138 -355 -131 -353
rect -138 -358 -133 -355
rect -112 -358 -104 -352
rect -102 -358 -97 -349
rect -95 -351 -88 -349
rect -95 -353 -92 -351
rect -90 -353 -88 -351
rect -95 -355 -88 -353
rect -95 -358 -90 -355
rect -241 -360 -235 -358
rect -241 -362 -239 -360
rect -237 -362 -235 -360
rect -241 -364 -235 -362
rect -198 -360 -192 -358
rect -198 -362 -196 -360
rect -194 -362 -192 -360
rect -198 -364 -192 -362
rect -155 -360 -149 -358
rect -155 -362 -153 -360
rect -151 -362 -149 -360
rect -155 -364 -149 -362
rect -112 -360 -106 -358
rect -112 -362 -110 -360
rect -108 -362 -106 -360
rect -112 -364 -106 -362
rect 267 146 274 148
rect 267 144 269 146
rect 271 144 274 146
rect 267 142 274 144
rect 276 145 284 148
rect 310 146 317 148
rect 276 142 286 145
rect 278 136 286 142
rect 288 136 293 145
rect 295 143 302 145
rect 295 141 298 143
rect 300 141 302 143
rect 310 144 312 146
rect 314 144 317 146
rect 310 142 317 144
rect 319 145 327 148
rect 353 146 360 148
rect 319 142 329 145
rect 295 139 302 141
rect 295 136 300 139
rect 321 136 329 142
rect 331 136 336 145
rect 338 143 345 145
rect 338 141 341 143
rect 343 141 345 143
rect 353 144 355 146
rect 357 144 360 146
rect 353 142 360 144
rect 362 145 370 148
rect 396 146 403 148
rect 362 142 372 145
rect 338 139 345 141
rect 338 136 343 139
rect 364 136 372 142
rect 374 136 379 145
rect 381 143 388 145
rect 381 141 384 143
rect 386 141 388 143
rect 396 144 398 146
rect 400 144 403 146
rect 396 142 403 144
rect 405 145 413 148
rect 405 142 415 145
rect 381 139 388 141
rect 381 136 386 139
rect 407 136 415 142
rect 417 136 422 145
rect 424 143 431 145
rect 424 141 427 143
rect 429 141 431 143
rect 424 139 431 141
rect 424 136 429 139
rect 278 134 284 136
rect 278 132 280 134
rect 282 132 284 134
rect 278 130 284 132
rect 321 134 327 136
rect 321 132 323 134
rect 325 132 327 134
rect 321 130 327 132
rect 364 134 370 136
rect 364 132 366 134
rect 368 132 370 134
rect 364 130 370 132
rect 407 134 413 136
rect 407 132 409 134
rect 411 132 413 134
rect 407 130 413 132
rect 288 50 293 57
rect 266 48 273 50
rect 266 46 268 48
rect 270 46 273 48
rect 266 44 273 46
rect 268 37 273 44
rect 275 44 283 50
rect 275 42 278 44
rect 280 42 283 44
rect 275 40 283 42
rect 285 47 293 50
rect 285 45 288 47
rect 290 45 293 47
rect 285 43 293 45
rect 295 55 303 57
rect 295 53 298 55
rect 300 53 303 55
rect 295 43 303 53
rect 305 55 312 57
rect 305 53 308 55
rect 310 53 312 55
rect 305 48 312 53
rect 318 50 323 57
rect 305 46 308 48
rect 310 46 312 48
rect 305 43 312 46
rect 316 48 323 50
rect 316 46 318 48
rect 320 46 323 48
rect 316 44 323 46
rect 285 40 290 43
rect 275 37 280 40
rect 318 37 323 44
rect 325 37 330 57
rect 332 51 339 57
rect 379 51 386 57
rect 332 41 341 51
rect 332 39 335 41
rect 337 39 341 41
rect 332 37 341 39
rect 343 48 350 51
rect 343 46 346 48
rect 348 46 350 48
rect 343 44 350 46
rect 368 48 375 51
rect 368 46 370 48
rect 372 46 375 48
rect 368 44 375 46
rect 343 37 348 44
rect 370 37 375 44
rect 377 41 386 51
rect 377 39 381 41
rect 383 39 386 41
rect 377 37 386 39
rect 388 37 393 57
rect 395 50 400 57
rect 406 55 413 57
rect 406 53 408 55
rect 410 53 413 55
rect 395 48 402 50
rect 395 46 398 48
rect 400 46 402 48
rect 395 44 402 46
rect 406 48 413 53
rect 406 46 408 48
rect 410 46 413 48
rect 395 37 400 44
rect 406 43 413 46
rect 415 55 423 57
rect 415 53 418 55
rect 420 53 423 55
rect 415 43 423 53
rect 425 50 430 57
rect 425 47 433 50
rect 425 45 428 47
rect 430 45 433 47
rect 425 43 433 45
rect 428 40 433 43
rect 435 44 443 50
rect 435 42 438 44
rect 440 42 443 44
rect 435 40 443 42
rect 438 37 443 40
rect 445 48 452 50
rect 445 46 448 48
rect 450 46 452 48
rect 445 44 452 46
rect 445 37 450 44
rect 28 -136 35 -130
rect 17 -139 24 -136
rect 17 -141 19 -139
rect 21 -141 24 -139
rect 17 -143 24 -141
rect 19 -150 24 -143
rect 26 -146 35 -136
rect 26 -148 30 -146
rect 32 -148 35 -146
rect 26 -150 35 -148
rect 37 -150 42 -130
rect 44 -137 49 -130
rect 55 -132 62 -130
rect 55 -134 57 -132
rect 59 -134 62 -132
rect 44 -139 51 -137
rect 44 -141 47 -139
rect 49 -141 51 -139
rect 44 -143 51 -141
rect 55 -139 62 -134
rect 55 -141 57 -139
rect 59 -141 62 -139
rect 44 -150 49 -143
rect 55 -144 62 -141
rect 64 -132 72 -130
rect 64 -134 67 -132
rect 69 -134 72 -132
rect 64 -144 72 -134
rect 74 -137 79 -130
rect 105 -137 112 -135
rect 74 -140 82 -137
rect 74 -142 77 -140
rect 79 -142 82 -140
rect 74 -144 82 -142
rect 77 -147 82 -144
rect 84 -143 92 -137
rect 84 -145 87 -143
rect 89 -145 92 -143
rect 84 -147 92 -145
rect 87 -150 92 -147
rect 94 -139 101 -137
rect 94 -141 97 -139
rect 99 -141 101 -139
rect 105 -139 107 -137
rect 109 -139 112 -137
rect 105 -141 112 -139
rect 114 -137 122 -135
rect 114 -139 117 -137
rect 119 -139 122 -137
rect 114 -141 122 -139
rect 124 -137 132 -135
rect 124 -139 127 -137
rect 129 -139 132 -137
rect 124 -141 132 -139
rect 134 -137 141 -135
rect 157 -136 164 -130
rect 134 -139 137 -137
rect 139 -139 141 -137
rect 134 -141 141 -139
rect 146 -139 153 -136
rect 146 -141 148 -139
rect 150 -141 153 -139
rect 94 -143 101 -141
rect 94 -150 99 -143
rect 146 -143 153 -141
rect 148 -150 153 -143
rect 155 -146 164 -136
rect 155 -148 159 -146
rect 161 -148 164 -146
rect 155 -150 164 -148
rect 166 -150 171 -130
rect 173 -137 178 -130
rect 184 -132 191 -130
rect 184 -134 186 -132
rect 188 -134 191 -132
rect 173 -139 180 -137
rect 173 -141 176 -139
rect 178 -141 180 -139
rect 173 -143 180 -141
rect 184 -139 191 -134
rect 184 -141 186 -139
rect 188 -141 191 -139
rect 173 -150 178 -143
rect 184 -144 191 -141
rect 193 -132 201 -130
rect 193 -134 196 -132
rect 198 -134 201 -132
rect 193 -144 201 -134
rect 203 -137 208 -130
rect 258 -137 263 -130
rect 203 -140 211 -137
rect 203 -142 206 -140
rect 208 -142 211 -140
rect 203 -144 211 -142
rect 206 -147 211 -144
rect 213 -143 221 -137
rect 213 -145 216 -143
rect 218 -145 221 -143
rect 213 -147 221 -145
rect 216 -150 221 -147
rect 223 -139 230 -137
rect 223 -141 226 -139
rect 228 -141 230 -139
rect 223 -143 230 -141
rect 236 -139 243 -137
rect 236 -141 238 -139
rect 240 -141 243 -139
rect 236 -143 243 -141
rect 223 -150 228 -143
rect 238 -150 243 -143
rect 245 -143 253 -137
rect 245 -145 248 -143
rect 250 -145 253 -143
rect 245 -147 253 -145
rect 255 -140 263 -137
rect 255 -142 258 -140
rect 260 -142 263 -140
rect 255 -144 263 -142
rect 265 -132 273 -130
rect 265 -134 268 -132
rect 270 -134 273 -132
rect 265 -144 273 -134
rect 275 -132 282 -130
rect 275 -134 278 -132
rect 280 -134 282 -132
rect 275 -139 282 -134
rect 288 -137 293 -130
rect 275 -141 278 -139
rect 280 -141 282 -139
rect 275 -144 282 -141
rect 286 -139 293 -137
rect 286 -141 288 -139
rect 290 -141 293 -139
rect 286 -143 293 -141
rect 255 -147 260 -144
rect 245 -150 250 -147
rect 288 -150 293 -143
rect 295 -150 300 -130
rect 302 -136 309 -130
rect 302 -146 311 -136
rect 302 -148 305 -146
rect 307 -148 311 -146
rect 302 -150 311 -148
rect 313 -139 320 -136
rect 313 -141 316 -139
rect 318 -141 320 -139
rect 325 -137 332 -135
rect 325 -139 327 -137
rect 329 -139 332 -137
rect 325 -141 332 -139
rect 334 -137 342 -135
rect 334 -139 337 -137
rect 339 -139 342 -137
rect 334 -141 342 -139
rect 344 -137 352 -135
rect 344 -139 347 -137
rect 349 -139 352 -137
rect 344 -141 352 -139
rect 354 -137 361 -135
rect 387 -137 392 -130
rect 354 -139 357 -137
rect 359 -139 361 -137
rect 354 -141 361 -139
rect 365 -139 372 -137
rect 365 -141 367 -139
rect 369 -141 372 -139
rect 313 -143 320 -141
rect 313 -150 318 -143
rect 365 -143 372 -141
rect 367 -150 372 -143
rect 374 -143 382 -137
rect 374 -145 377 -143
rect 379 -145 382 -143
rect 374 -147 382 -145
rect 384 -140 392 -137
rect 384 -142 387 -140
rect 389 -142 392 -140
rect 384 -144 392 -142
rect 394 -132 402 -130
rect 394 -134 397 -132
rect 399 -134 402 -132
rect 394 -144 402 -134
rect 404 -132 411 -130
rect 404 -134 407 -132
rect 409 -134 411 -132
rect 404 -139 411 -134
rect 417 -137 422 -130
rect 404 -141 407 -139
rect 409 -141 411 -139
rect 404 -144 411 -141
rect 415 -139 422 -137
rect 415 -141 417 -139
rect 419 -141 422 -139
rect 415 -143 422 -141
rect 384 -147 389 -144
rect 374 -150 379 -147
rect 417 -150 422 -143
rect 424 -150 429 -130
rect 431 -136 438 -130
rect 466 -136 473 -130
rect 431 -146 440 -136
rect 431 -148 434 -146
rect 436 -148 440 -146
rect 431 -150 440 -148
rect 442 -139 449 -136
rect 442 -141 445 -139
rect 447 -141 449 -139
rect 442 -143 449 -141
rect 455 -139 462 -136
rect 455 -141 457 -139
rect 459 -141 462 -139
rect 455 -143 462 -141
rect 442 -150 447 -143
rect 457 -150 462 -143
rect 464 -146 473 -136
rect 464 -148 468 -146
rect 470 -148 473 -146
rect 464 -150 473 -148
rect 475 -150 480 -130
rect 482 -137 487 -130
rect 493 -132 500 -130
rect 493 -134 495 -132
rect 497 -134 500 -132
rect 482 -139 489 -137
rect 482 -141 485 -139
rect 487 -141 489 -139
rect 482 -143 489 -141
rect 493 -139 500 -134
rect 493 -141 495 -139
rect 497 -141 500 -139
rect 482 -150 487 -143
rect 493 -144 500 -141
rect 502 -132 510 -130
rect 502 -134 505 -132
rect 507 -134 510 -132
rect 502 -144 510 -134
rect 512 -137 517 -130
rect 543 -137 550 -135
rect 512 -140 520 -137
rect 512 -142 515 -140
rect 517 -142 520 -140
rect 512 -144 520 -142
rect 515 -147 520 -144
rect 522 -143 530 -137
rect 522 -145 525 -143
rect 527 -145 530 -143
rect 522 -147 530 -145
rect 525 -150 530 -147
rect 532 -139 539 -137
rect 532 -141 535 -139
rect 537 -141 539 -139
rect 543 -139 545 -137
rect 547 -139 550 -137
rect 543 -141 550 -139
rect 552 -137 560 -135
rect 552 -139 555 -137
rect 557 -139 560 -137
rect 552 -141 560 -139
rect 562 -137 570 -135
rect 562 -139 565 -137
rect 567 -139 570 -137
rect 562 -141 570 -139
rect 572 -137 579 -135
rect 595 -136 602 -130
rect 572 -139 575 -137
rect 577 -139 579 -137
rect 572 -141 579 -139
rect 584 -139 591 -136
rect 584 -141 586 -139
rect 588 -141 591 -139
rect 532 -143 539 -141
rect 532 -150 537 -143
rect 584 -143 591 -141
rect 586 -150 591 -143
rect 593 -146 602 -136
rect 593 -148 597 -146
rect 599 -148 602 -146
rect 593 -150 602 -148
rect 604 -150 609 -130
rect 611 -137 616 -130
rect 622 -132 629 -130
rect 622 -134 624 -132
rect 626 -134 629 -132
rect 611 -139 618 -137
rect 611 -141 614 -139
rect 616 -141 618 -139
rect 611 -143 618 -141
rect 622 -139 629 -134
rect 622 -141 624 -139
rect 626 -141 629 -139
rect 611 -150 616 -143
rect 622 -144 629 -141
rect 631 -132 639 -130
rect 631 -134 634 -132
rect 636 -134 639 -132
rect 631 -144 639 -134
rect 641 -137 646 -130
rect 687 -136 694 -130
rect 641 -140 649 -137
rect 641 -142 644 -140
rect 646 -142 649 -140
rect 641 -144 649 -142
rect 644 -147 649 -144
rect 651 -143 659 -137
rect 651 -145 654 -143
rect 656 -145 659 -143
rect 651 -147 659 -145
rect 654 -150 659 -147
rect 661 -139 668 -137
rect 661 -141 664 -139
rect 666 -141 668 -139
rect 661 -143 668 -141
rect 676 -139 683 -136
rect 676 -141 678 -139
rect 680 -141 683 -139
rect 676 -143 683 -141
rect 661 -150 666 -143
rect 678 -150 683 -143
rect 685 -146 694 -136
rect 685 -148 689 -146
rect 691 -148 694 -146
rect 685 -150 694 -148
rect 696 -150 701 -130
rect 703 -137 708 -130
rect 714 -132 721 -130
rect 714 -134 716 -132
rect 718 -134 721 -132
rect 703 -139 710 -137
rect 703 -141 706 -139
rect 708 -141 710 -139
rect 703 -143 710 -141
rect 714 -139 721 -134
rect 714 -141 716 -139
rect 718 -141 721 -139
rect 703 -150 708 -143
rect 714 -144 721 -141
rect 723 -132 731 -130
rect 723 -134 726 -132
rect 728 -134 731 -132
rect 723 -144 731 -134
rect 733 -137 738 -130
rect 733 -140 741 -137
rect 733 -142 736 -140
rect 738 -142 741 -140
rect 733 -144 741 -142
rect 736 -147 741 -144
rect 743 -143 751 -137
rect 743 -145 746 -143
rect 748 -145 751 -143
rect 743 -147 751 -145
rect 746 -150 751 -147
rect 753 -139 760 -137
rect 753 -141 756 -139
rect 758 -141 760 -139
rect 753 -143 760 -141
rect 753 -150 758 -143
rect 400 -271 407 -269
rect 400 -273 402 -271
rect 404 -273 407 -271
rect 400 -275 407 -273
rect 409 -272 417 -269
rect 443 -271 450 -269
rect 409 -275 419 -272
rect 411 -281 419 -275
rect 421 -281 426 -272
rect 428 -274 435 -272
rect 428 -276 431 -274
rect 433 -276 435 -274
rect 443 -273 445 -271
rect 447 -273 450 -271
rect 443 -275 450 -273
rect 452 -272 460 -269
rect 486 -271 493 -269
rect 452 -275 462 -272
rect 428 -278 435 -276
rect 428 -281 433 -278
rect 454 -281 462 -275
rect 464 -281 469 -272
rect 471 -274 478 -272
rect 471 -276 474 -274
rect 476 -276 478 -274
rect 486 -273 488 -271
rect 490 -273 493 -271
rect 486 -275 493 -273
rect 495 -272 503 -269
rect 529 -271 536 -269
rect 495 -275 505 -272
rect 471 -278 478 -276
rect 471 -281 476 -278
rect 497 -281 505 -275
rect 507 -281 512 -272
rect 514 -274 521 -272
rect 514 -276 517 -274
rect 519 -276 521 -274
rect 529 -273 531 -271
rect 533 -273 536 -271
rect 529 -275 536 -273
rect 538 -272 546 -269
rect 538 -275 548 -272
rect 514 -278 521 -276
rect 514 -281 519 -278
rect 540 -281 548 -275
rect 550 -281 555 -272
rect 557 -274 564 -272
rect 557 -276 560 -274
rect 562 -276 564 -274
rect 557 -278 564 -276
rect 557 -281 562 -278
rect 411 -283 417 -281
rect 411 -285 413 -283
rect 415 -285 417 -283
rect 411 -287 417 -285
rect 454 -283 460 -281
rect 454 -285 456 -283
rect 458 -285 460 -283
rect 454 -287 460 -285
rect 497 -283 503 -281
rect 497 -285 499 -283
rect 501 -285 503 -283
rect 497 -287 503 -285
rect 540 -283 546 -281
rect 540 -285 542 -283
rect 544 -285 546 -283
rect 540 -287 546 -285
rect 421 -367 426 -360
rect 399 -369 406 -367
rect 399 -371 401 -369
rect 403 -371 406 -369
rect 399 -373 406 -371
rect 401 -380 406 -373
rect 408 -373 416 -367
rect 408 -375 411 -373
rect 413 -375 416 -373
rect 408 -377 416 -375
rect 418 -370 426 -367
rect 418 -372 421 -370
rect 423 -372 426 -370
rect 418 -374 426 -372
rect 428 -362 436 -360
rect 428 -364 431 -362
rect 433 -364 436 -362
rect 428 -374 436 -364
rect 438 -362 445 -360
rect 438 -364 441 -362
rect 443 -364 445 -362
rect 438 -369 445 -364
rect 451 -367 456 -360
rect 438 -371 441 -369
rect 443 -371 445 -369
rect 438 -374 445 -371
rect 449 -369 456 -367
rect 449 -371 451 -369
rect 453 -371 456 -369
rect 449 -373 456 -371
rect 418 -377 423 -374
rect 408 -380 413 -377
rect 451 -380 456 -373
rect 458 -380 463 -360
rect 465 -366 472 -360
rect 512 -366 519 -360
rect 465 -376 474 -366
rect 465 -378 468 -376
rect 470 -378 474 -376
rect 465 -380 474 -378
rect 476 -369 483 -366
rect 476 -371 479 -369
rect 481 -371 483 -369
rect 476 -373 483 -371
rect 501 -369 508 -366
rect 501 -371 503 -369
rect 505 -371 508 -369
rect 501 -373 508 -371
rect 476 -380 481 -373
rect 503 -380 508 -373
rect 510 -376 519 -366
rect 510 -378 514 -376
rect 516 -378 519 -376
rect 510 -380 519 -378
rect 521 -380 526 -360
rect 528 -367 533 -360
rect 539 -362 546 -360
rect 539 -364 541 -362
rect 543 -364 546 -362
rect 528 -369 535 -367
rect 528 -371 531 -369
rect 533 -371 535 -369
rect 528 -373 535 -371
rect 539 -369 546 -364
rect 539 -371 541 -369
rect 543 -371 546 -369
rect 528 -380 533 -373
rect 539 -374 546 -371
rect 548 -362 556 -360
rect 548 -364 551 -362
rect 553 -364 556 -362
rect 548 -374 556 -364
rect 558 -367 563 -360
rect 558 -370 566 -367
rect 558 -372 561 -370
rect 563 -372 566 -370
rect 558 -374 566 -372
rect 561 -377 566 -374
rect 568 -373 576 -367
rect 568 -375 571 -373
rect 573 -375 576 -373
rect 568 -377 576 -375
rect 571 -380 576 -377
rect 578 -369 585 -367
rect 578 -371 581 -369
rect 583 -371 585 -369
rect 578 -373 585 -371
rect 578 -380 583 -373
rect -231 -444 -226 -437
rect -253 -446 -246 -444
rect -253 -448 -251 -446
rect -249 -448 -246 -446
rect -253 -450 -246 -448
rect -251 -457 -246 -450
rect -244 -450 -236 -444
rect -244 -452 -241 -450
rect -239 -452 -236 -450
rect -244 -454 -236 -452
rect -234 -447 -226 -444
rect -234 -449 -231 -447
rect -229 -449 -226 -447
rect -234 -451 -226 -449
rect -224 -439 -216 -437
rect -224 -441 -221 -439
rect -219 -441 -216 -439
rect -224 -451 -216 -441
rect -214 -439 -207 -437
rect -214 -441 -211 -439
rect -209 -441 -207 -439
rect -214 -446 -207 -441
rect -201 -444 -196 -437
rect -214 -448 -211 -446
rect -209 -448 -207 -446
rect -214 -451 -207 -448
rect -203 -446 -196 -444
rect -203 -448 -201 -446
rect -199 -448 -196 -446
rect -203 -450 -196 -448
rect -234 -454 -229 -451
rect -244 -457 -239 -454
rect -201 -457 -196 -450
rect -194 -457 -189 -437
rect -187 -443 -180 -437
rect -140 -443 -133 -437
rect -187 -453 -178 -443
rect -187 -455 -184 -453
rect -182 -455 -178 -453
rect -187 -457 -178 -455
rect -176 -446 -169 -443
rect -176 -448 -173 -446
rect -171 -448 -169 -446
rect -176 -450 -169 -448
rect -151 -446 -144 -443
rect -151 -448 -149 -446
rect -147 -448 -144 -446
rect -151 -450 -144 -448
rect -176 -457 -171 -450
rect -149 -457 -144 -450
rect -142 -453 -133 -443
rect -142 -455 -138 -453
rect -136 -455 -133 -453
rect -142 -457 -133 -455
rect -131 -457 -126 -437
rect -124 -444 -119 -437
rect -113 -439 -106 -437
rect -113 -441 -111 -439
rect -109 -441 -106 -439
rect -124 -446 -117 -444
rect -124 -448 -121 -446
rect -119 -448 -117 -446
rect -124 -450 -117 -448
rect -113 -446 -106 -441
rect -113 -448 -111 -446
rect -109 -448 -106 -446
rect -124 -457 -119 -450
rect -113 -451 -106 -448
rect -104 -439 -96 -437
rect -104 -441 -101 -439
rect -99 -441 -96 -439
rect -104 -451 -96 -441
rect -94 -444 -89 -437
rect -94 -447 -86 -444
rect -94 -449 -91 -447
rect -89 -449 -86 -447
rect -94 -451 -86 -449
rect -91 -454 -86 -451
rect -84 -450 -76 -444
rect -84 -452 -81 -450
rect -79 -452 -76 -450
rect -84 -454 -76 -452
rect -81 -457 -76 -454
rect -74 -446 -67 -444
rect -74 -448 -71 -446
rect -69 -448 -67 -446
rect -74 -450 -67 -448
rect -74 -457 -69 -450
rect 30 -521 37 -515
rect 19 -524 26 -521
rect 19 -526 21 -524
rect 23 -526 26 -524
rect 19 -528 26 -526
rect 21 -535 26 -528
rect 28 -531 37 -521
rect 28 -533 32 -531
rect 34 -533 37 -531
rect 28 -535 37 -533
rect 39 -535 44 -515
rect 46 -522 51 -515
rect 57 -517 64 -515
rect 57 -519 59 -517
rect 61 -519 64 -517
rect 46 -524 53 -522
rect 46 -526 49 -524
rect 51 -526 53 -524
rect 46 -528 53 -526
rect 57 -524 64 -519
rect 57 -526 59 -524
rect 61 -526 64 -524
rect 46 -535 51 -528
rect 57 -529 64 -526
rect 66 -517 74 -515
rect 66 -519 69 -517
rect 71 -519 74 -517
rect 66 -529 74 -519
rect 76 -522 81 -515
rect 107 -522 114 -520
rect 76 -525 84 -522
rect 76 -527 79 -525
rect 81 -527 84 -525
rect 76 -529 84 -527
rect 79 -532 84 -529
rect 86 -528 94 -522
rect 86 -530 89 -528
rect 91 -530 94 -528
rect 86 -532 94 -530
rect 89 -535 94 -532
rect 96 -524 103 -522
rect 96 -526 99 -524
rect 101 -526 103 -524
rect 107 -524 109 -522
rect 111 -524 114 -522
rect 107 -526 114 -524
rect 116 -522 124 -520
rect 116 -524 119 -522
rect 121 -524 124 -522
rect 116 -526 124 -524
rect 126 -522 134 -520
rect 126 -524 129 -522
rect 131 -524 134 -522
rect 126 -526 134 -524
rect 136 -522 143 -520
rect 159 -521 166 -515
rect 136 -524 139 -522
rect 141 -524 143 -522
rect 136 -526 143 -524
rect 148 -524 155 -521
rect 148 -526 150 -524
rect 152 -526 155 -524
rect 96 -528 103 -526
rect 96 -535 101 -528
rect 148 -528 155 -526
rect 150 -535 155 -528
rect 157 -531 166 -521
rect 157 -533 161 -531
rect 163 -533 166 -531
rect 157 -535 166 -533
rect 168 -535 173 -515
rect 175 -522 180 -515
rect 186 -517 193 -515
rect 186 -519 188 -517
rect 190 -519 193 -517
rect 175 -524 182 -522
rect 175 -526 178 -524
rect 180 -526 182 -524
rect 175 -528 182 -526
rect 186 -524 193 -519
rect 186 -526 188 -524
rect 190 -526 193 -524
rect 175 -535 180 -528
rect 186 -529 193 -526
rect 195 -517 203 -515
rect 195 -519 198 -517
rect 200 -519 203 -517
rect 195 -529 203 -519
rect 205 -522 210 -515
rect 260 -522 265 -515
rect 205 -525 213 -522
rect 205 -527 208 -525
rect 210 -527 213 -525
rect 205 -529 213 -527
rect 208 -532 213 -529
rect 215 -528 223 -522
rect 215 -530 218 -528
rect 220 -530 223 -528
rect 215 -532 223 -530
rect 218 -535 223 -532
rect 225 -524 232 -522
rect 225 -526 228 -524
rect 230 -526 232 -524
rect 225 -528 232 -526
rect 238 -524 245 -522
rect 238 -526 240 -524
rect 242 -526 245 -524
rect 238 -528 245 -526
rect 225 -535 230 -528
rect 240 -535 245 -528
rect 247 -528 255 -522
rect 247 -530 250 -528
rect 252 -530 255 -528
rect 247 -532 255 -530
rect 257 -525 265 -522
rect 257 -527 260 -525
rect 262 -527 265 -525
rect 257 -529 265 -527
rect 267 -517 275 -515
rect 267 -519 270 -517
rect 272 -519 275 -517
rect 267 -529 275 -519
rect 277 -517 284 -515
rect 277 -519 280 -517
rect 282 -519 284 -517
rect 277 -524 284 -519
rect 290 -522 295 -515
rect 277 -526 280 -524
rect 282 -526 284 -524
rect 277 -529 284 -526
rect 288 -524 295 -522
rect 288 -526 290 -524
rect 292 -526 295 -524
rect 288 -528 295 -526
rect 257 -532 262 -529
rect 247 -535 252 -532
rect 290 -535 295 -528
rect 297 -535 302 -515
rect 304 -521 311 -515
rect 304 -531 313 -521
rect 304 -533 307 -531
rect 309 -533 313 -531
rect 304 -535 313 -533
rect 315 -524 322 -521
rect 315 -526 318 -524
rect 320 -526 322 -524
rect 327 -522 334 -520
rect 327 -524 329 -522
rect 331 -524 334 -522
rect 327 -526 334 -524
rect 336 -522 344 -520
rect 336 -524 339 -522
rect 341 -524 344 -522
rect 336 -526 344 -524
rect 346 -522 354 -520
rect 346 -524 349 -522
rect 351 -524 354 -522
rect 346 -526 354 -524
rect 356 -522 363 -520
rect 389 -522 394 -515
rect 356 -524 359 -522
rect 361 -524 363 -522
rect 356 -526 363 -524
rect 367 -524 374 -522
rect 367 -526 369 -524
rect 371 -526 374 -524
rect 315 -528 322 -526
rect 315 -535 320 -528
rect 367 -528 374 -526
rect 369 -535 374 -528
rect 376 -528 384 -522
rect 376 -530 379 -528
rect 381 -530 384 -528
rect 376 -532 384 -530
rect 386 -525 394 -522
rect 386 -527 389 -525
rect 391 -527 394 -525
rect 386 -529 394 -527
rect 396 -517 404 -515
rect 396 -519 399 -517
rect 401 -519 404 -517
rect 396 -529 404 -519
rect 406 -517 413 -515
rect 406 -519 409 -517
rect 411 -519 413 -517
rect 406 -524 413 -519
rect 419 -522 424 -515
rect 406 -526 409 -524
rect 411 -526 413 -524
rect 406 -529 413 -526
rect 417 -524 424 -522
rect 417 -526 419 -524
rect 421 -526 424 -524
rect 417 -528 424 -526
rect 386 -532 391 -529
rect 376 -535 381 -532
rect 419 -535 424 -528
rect 426 -535 431 -515
rect 433 -521 440 -515
rect 468 -521 475 -515
rect 433 -531 442 -521
rect 433 -533 436 -531
rect 438 -533 442 -531
rect 433 -535 442 -533
rect 444 -524 451 -521
rect 444 -526 447 -524
rect 449 -526 451 -524
rect 444 -528 451 -526
rect 457 -524 464 -521
rect 457 -526 459 -524
rect 461 -526 464 -524
rect 457 -528 464 -526
rect 444 -535 449 -528
rect 459 -535 464 -528
rect 466 -531 475 -521
rect 466 -533 470 -531
rect 472 -533 475 -531
rect 466 -535 475 -533
rect 477 -535 482 -515
rect 484 -522 489 -515
rect 495 -517 502 -515
rect 495 -519 497 -517
rect 499 -519 502 -517
rect 484 -524 491 -522
rect 484 -526 487 -524
rect 489 -526 491 -524
rect 484 -528 491 -526
rect 495 -524 502 -519
rect 495 -526 497 -524
rect 499 -526 502 -524
rect 484 -535 489 -528
rect 495 -529 502 -526
rect 504 -517 512 -515
rect 504 -519 507 -517
rect 509 -519 512 -517
rect 504 -529 512 -519
rect 514 -522 519 -515
rect 545 -522 552 -520
rect 514 -525 522 -522
rect 514 -527 517 -525
rect 519 -527 522 -525
rect 514 -529 522 -527
rect 517 -532 522 -529
rect 524 -528 532 -522
rect 524 -530 527 -528
rect 529 -530 532 -528
rect 524 -532 532 -530
rect 527 -535 532 -532
rect 534 -524 541 -522
rect 534 -526 537 -524
rect 539 -526 541 -524
rect 545 -524 547 -522
rect 549 -524 552 -522
rect 545 -526 552 -524
rect 554 -522 562 -520
rect 554 -524 557 -522
rect 559 -524 562 -522
rect 554 -526 562 -524
rect 564 -522 572 -520
rect 564 -524 567 -522
rect 569 -524 572 -522
rect 564 -526 572 -524
rect 574 -522 581 -520
rect 597 -521 604 -515
rect 574 -524 577 -522
rect 579 -524 581 -522
rect 574 -526 581 -524
rect 586 -524 593 -521
rect 586 -526 588 -524
rect 590 -526 593 -524
rect 534 -528 541 -526
rect 534 -535 539 -528
rect 586 -528 593 -526
rect 588 -535 593 -528
rect 595 -531 604 -521
rect 595 -533 599 -531
rect 601 -533 604 -531
rect 595 -535 604 -533
rect 606 -535 611 -515
rect 613 -522 618 -515
rect 624 -517 631 -515
rect 624 -519 626 -517
rect 628 -519 631 -517
rect 613 -524 620 -522
rect 613 -526 616 -524
rect 618 -526 620 -524
rect 613 -528 620 -526
rect 624 -524 631 -519
rect 624 -526 626 -524
rect 628 -526 631 -524
rect 613 -535 618 -528
rect 624 -529 631 -526
rect 633 -517 641 -515
rect 633 -519 636 -517
rect 638 -519 641 -517
rect 633 -529 641 -519
rect 643 -522 648 -515
rect 689 -521 696 -515
rect 643 -525 651 -522
rect 643 -527 646 -525
rect 648 -527 651 -525
rect 643 -529 651 -527
rect 646 -532 651 -529
rect 653 -528 661 -522
rect 653 -530 656 -528
rect 658 -530 661 -528
rect 653 -532 661 -530
rect 656 -535 661 -532
rect 663 -524 670 -522
rect 663 -526 666 -524
rect 668 -526 670 -524
rect 663 -528 670 -526
rect 678 -524 685 -521
rect 678 -526 680 -524
rect 682 -526 685 -524
rect 678 -528 685 -526
rect 663 -535 668 -528
rect 680 -535 685 -528
rect 687 -531 696 -521
rect 687 -533 691 -531
rect 693 -533 696 -531
rect 687 -535 696 -533
rect 698 -535 703 -515
rect 705 -522 710 -515
rect 716 -517 723 -515
rect 716 -519 718 -517
rect 720 -519 723 -517
rect 705 -524 712 -522
rect 705 -526 708 -524
rect 710 -526 712 -524
rect 705 -528 712 -526
rect 716 -524 723 -519
rect 716 -526 718 -524
rect 720 -526 723 -524
rect 705 -535 710 -528
rect 716 -529 723 -526
rect 725 -517 733 -515
rect 725 -519 728 -517
rect 730 -519 733 -517
rect 725 -529 733 -519
rect 735 -522 740 -515
rect 735 -525 743 -522
rect 735 -527 738 -525
rect 740 -527 743 -525
rect 735 -529 743 -527
rect 738 -532 743 -529
rect 745 -528 753 -522
rect 745 -530 748 -528
rect 750 -530 753 -528
rect 745 -532 753 -530
rect 748 -535 753 -532
rect 755 -524 762 -522
rect 755 -526 758 -524
rect 760 -526 762 -524
rect 755 -528 762 -526
rect 755 -535 760 -528
rect -237 -655 -230 -649
rect -248 -658 -241 -655
rect -248 -660 -246 -658
rect -244 -660 -241 -658
rect -248 -662 -241 -660
rect -246 -669 -241 -662
rect -239 -665 -230 -655
rect -239 -667 -235 -665
rect -233 -667 -230 -665
rect -239 -669 -230 -667
rect -228 -669 -223 -649
rect -221 -656 -216 -649
rect -210 -651 -203 -649
rect -210 -653 -208 -651
rect -206 -653 -203 -651
rect -221 -658 -214 -656
rect -221 -660 -218 -658
rect -216 -660 -214 -658
rect -221 -662 -214 -660
rect -210 -658 -203 -653
rect -210 -660 -208 -658
rect -206 -660 -203 -658
rect -221 -669 -216 -662
rect -210 -663 -203 -660
rect -201 -651 -193 -649
rect -201 -653 -198 -651
rect -196 -653 -193 -651
rect -201 -663 -193 -653
rect -191 -656 -186 -649
rect -160 -656 -153 -654
rect -191 -659 -183 -656
rect -191 -661 -188 -659
rect -186 -661 -183 -659
rect -191 -663 -183 -661
rect -188 -666 -183 -663
rect -181 -662 -173 -656
rect -181 -664 -178 -662
rect -176 -664 -173 -662
rect -181 -666 -173 -664
rect -178 -669 -173 -666
rect -171 -658 -164 -656
rect -171 -660 -168 -658
rect -166 -660 -164 -658
rect -160 -658 -158 -656
rect -156 -658 -153 -656
rect -160 -660 -153 -658
rect -151 -656 -143 -654
rect -151 -658 -148 -656
rect -146 -658 -143 -656
rect -151 -660 -143 -658
rect -141 -656 -133 -654
rect -141 -658 -138 -656
rect -136 -658 -133 -656
rect -141 -660 -133 -658
rect -131 -656 -124 -654
rect -108 -655 -101 -649
rect -131 -658 -128 -656
rect -126 -658 -124 -656
rect -131 -660 -124 -658
rect -119 -658 -112 -655
rect -119 -660 -117 -658
rect -115 -660 -112 -658
rect -171 -662 -164 -660
rect -171 -669 -166 -662
rect -119 -662 -112 -660
rect -117 -669 -112 -662
rect -110 -665 -101 -655
rect -110 -667 -106 -665
rect -104 -667 -101 -665
rect -110 -669 -101 -667
rect -99 -669 -94 -649
rect -92 -656 -87 -649
rect -81 -651 -74 -649
rect -81 -653 -79 -651
rect -77 -653 -74 -651
rect -92 -658 -85 -656
rect -92 -660 -89 -658
rect -87 -660 -85 -658
rect -92 -662 -85 -660
rect -81 -658 -74 -653
rect -81 -660 -79 -658
rect -77 -660 -74 -658
rect -92 -669 -87 -662
rect -81 -663 -74 -660
rect -72 -651 -64 -649
rect -72 -653 -69 -651
rect -67 -653 -64 -651
rect -72 -663 -64 -653
rect -62 -656 -57 -649
rect -7 -656 -2 -649
rect -62 -659 -54 -656
rect -62 -661 -59 -659
rect -57 -661 -54 -659
rect -62 -663 -54 -661
rect -59 -666 -54 -663
rect -52 -662 -44 -656
rect -52 -664 -49 -662
rect -47 -664 -44 -662
rect -52 -666 -44 -664
rect -49 -669 -44 -666
rect -42 -658 -35 -656
rect -42 -660 -39 -658
rect -37 -660 -35 -658
rect -42 -662 -35 -660
rect -29 -658 -22 -656
rect -29 -660 -27 -658
rect -25 -660 -22 -658
rect -29 -662 -22 -660
rect -42 -669 -37 -662
rect -27 -669 -22 -662
rect -20 -662 -12 -656
rect -20 -664 -17 -662
rect -15 -664 -12 -662
rect -20 -666 -12 -664
rect -10 -659 -2 -656
rect -10 -661 -7 -659
rect -5 -661 -2 -659
rect -10 -663 -2 -661
rect 0 -651 8 -649
rect 0 -653 3 -651
rect 5 -653 8 -651
rect 0 -663 8 -653
rect 10 -651 17 -649
rect 10 -653 13 -651
rect 15 -653 17 -651
rect 10 -658 17 -653
rect 23 -656 28 -649
rect 10 -660 13 -658
rect 15 -660 17 -658
rect 10 -663 17 -660
rect 21 -658 28 -656
rect 21 -660 23 -658
rect 25 -660 28 -658
rect 21 -662 28 -660
rect -10 -666 -5 -663
rect -20 -669 -15 -666
rect 23 -669 28 -662
rect 30 -669 35 -649
rect 37 -655 44 -649
rect 37 -665 46 -655
rect 37 -667 40 -665
rect 42 -667 46 -665
rect 37 -669 46 -667
rect 48 -658 55 -655
rect 48 -660 51 -658
rect 53 -660 55 -658
rect 60 -656 67 -654
rect 60 -658 62 -656
rect 64 -658 67 -656
rect 60 -660 67 -658
rect 69 -656 77 -654
rect 69 -658 72 -656
rect 74 -658 77 -656
rect 69 -660 77 -658
rect 79 -656 87 -654
rect 79 -658 82 -656
rect 84 -658 87 -656
rect 79 -660 87 -658
rect 89 -656 96 -654
rect 122 -656 127 -649
rect 89 -658 92 -656
rect 94 -658 96 -656
rect 89 -660 96 -658
rect 100 -658 107 -656
rect 100 -660 102 -658
rect 104 -660 107 -658
rect 48 -662 55 -660
rect 48 -669 53 -662
rect 100 -662 107 -660
rect 102 -669 107 -662
rect 109 -662 117 -656
rect 109 -664 112 -662
rect 114 -664 117 -662
rect 109 -666 117 -664
rect 119 -659 127 -656
rect 119 -661 122 -659
rect 124 -661 127 -659
rect 119 -663 127 -661
rect 129 -651 137 -649
rect 129 -653 132 -651
rect 134 -653 137 -651
rect 129 -663 137 -653
rect 139 -651 146 -649
rect 139 -653 142 -651
rect 144 -653 146 -651
rect 139 -658 146 -653
rect 152 -656 157 -649
rect 139 -660 142 -658
rect 144 -660 146 -658
rect 139 -663 146 -660
rect 150 -658 157 -656
rect 150 -660 152 -658
rect 154 -660 157 -658
rect 150 -662 157 -660
rect 119 -666 124 -663
rect 109 -669 114 -666
rect 152 -669 157 -662
rect 159 -669 164 -649
rect 166 -655 173 -649
rect 201 -655 208 -649
rect 166 -665 175 -655
rect 166 -667 169 -665
rect 171 -667 175 -665
rect 166 -669 175 -667
rect 177 -658 184 -655
rect 177 -660 180 -658
rect 182 -660 184 -658
rect 177 -662 184 -660
rect 190 -658 197 -655
rect 190 -660 192 -658
rect 194 -660 197 -658
rect 190 -662 197 -660
rect 177 -669 182 -662
rect 192 -669 197 -662
rect 199 -665 208 -655
rect 199 -667 203 -665
rect 205 -667 208 -665
rect 199 -669 208 -667
rect 210 -669 215 -649
rect 217 -656 222 -649
rect 228 -651 235 -649
rect 228 -653 230 -651
rect 232 -653 235 -651
rect 217 -658 224 -656
rect 217 -660 220 -658
rect 222 -660 224 -658
rect 217 -662 224 -660
rect 228 -658 235 -653
rect 228 -660 230 -658
rect 232 -660 235 -658
rect 217 -669 222 -662
rect 228 -663 235 -660
rect 237 -651 245 -649
rect 237 -653 240 -651
rect 242 -653 245 -651
rect 237 -663 245 -653
rect 247 -656 252 -649
rect 278 -656 285 -654
rect 247 -659 255 -656
rect 247 -661 250 -659
rect 252 -661 255 -659
rect 247 -663 255 -661
rect 250 -666 255 -663
rect 257 -662 265 -656
rect 257 -664 260 -662
rect 262 -664 265 -662
rect 257 -666 265 -664
rect 260 -669 265 -666
rect 267 -658 274 -656
rect 267 -660 270 -658
rect 272 -660 274 -658
rect 278 -658 280 -656
rect 282 -658 285 -656
rect 278 -660 285 -658
rect 287 -656 295 -654
rect 287 -658 290 -656
rect 292 -658 295 -656
rect 287 -660 295 -658
rect 297 -656 305 -654
rect 297 -658 300 -656
rect 302 -658 305 -656
rect 297 -660 305 -658
rect 307 -656 314 -654
rect 330 -655 337 -649
rect 307 -658 310 -656
rect 312 -658 314 -656
rect 307 -660 314 -658
rect 319 -658 326 -655
rect 319 -660 321 -658
rect 323 -660 326 -658
rect 267 -662 274 -660
rect 267 -669 272 -662
rect 319 -662 326 -660
rect 321 -669 326 -662
rect 328 -665 337 -655
rect 328 -667 332 -665
rect 334 -667 337 -665
rect 328 -669 337 -667
rect 339 -669 344 -649
rect 346 -656 351 -649
rect 357 -651 364 -649
rect 357 -653 359 -651
rect 361 -653 364 -651
rect 346 -658 353 -656
rect 346 -660 349 -658
rect 351 -660 353 -658
rect 346 -662 353 -660
rect 357 -658 364 -653
rect 357 -660 359 -658
rect 361 -660 364 -658
rect 346 -669 351 -662
rect 357 -663 364 -660
rect 366 -651 374 -649
rect 366 -653 369 -651
rect 371 -653 374 -651
rect 366 -663 374 -653
rect 376 -656 381 -649
rect 422 -655 429 -649
rect 376 -659 384 -656
rect 376 -661 379 -659
rect 381 -661 384 -659
rect 376 -663 384 -661
rect 379 -666 384 -663
rect 386 -662 394 -656
rect 386 -664 389 -662
rect 391 -664 394 -662
rect 386 -666 394 -664
rect 389 -669 394 -666
rect 396 -658 403 -656
rect 396 -660 399 -658
rect 401 -660 403 -658
rect 396 -662 403 -660
rect 411 -658 418 -655
rect 411 -660 413 -658
rect 415 -660 418 -658
rect 411 -662 418 -660
rect 396 -669 401 -662
rect 413 -669 418 -662
rect 420 -665 429 -655
rect 420 -667 424 -665
rect 426 -667 429 -665
rect 420 -669 429 -667
rect 431 -669 436 -649
rect 438 -656 443 -649
rect 449 -651 456 -649
rect 449 -653 451 -651
rect 453 -653 456 -651
rect 438 -658 445 -656
rect 438 -660 441 -658
rect 443 -660 445 -658
rect 438 -662 445 -660
rect 449 -658 456 -653
rect 449 -660 451 -658
rect 453 -660 456 -658
rect 438 -669 443 -662
rect 449 -663 456 -660
rect 458 -651 466 -649
rect 458 -653 461 -651
rect 463 -653 466 -651
rect 458 -663 466 -653
rect 468 -656 473 -649
rect 468 -659 476 -656
rect 468 -661 471 -659
rect 473 -661 476 -659
rect 468 -663 476 -661
rect 471 -666 476 -663
rect 478 -662 486 -656
rect 478 -664 481 -662
rect 483 -664 486 -662
rect 478 -666 486 -664
rect 481 -669 486 -666
rect 488 -658 495 -656
rect 488 -660 491 -658
rect 493 -660 495 -658
rect 488 -662 495 -660
rect 488 -669 493 -662
<< pdif >>
rect -251 -71 -246 -65
rect -253 -73 -246 -71
rect -253 -75 -251 -73
rect -249 -75 -246 -73
rect -253 -77 -246 -75
rect -244 -67 -238 -65
rect -244 -73 -236 -67
rect -244 -75 -241 -73
rect -239 -75 -236 -73
rect -244 -77 -236 -75
rect -234 -73 -226 -67
rect -234 -75 -231 -73
rect -229 -75 -226 -73
rect -234 -77 -226 -75
rect -224 -69 -217 -67
rect -224 -71 -221 -69
rect -219 -71 -217 -69
rect -208 -71 -203 -65
rect -224 -77 -217 -71
rect -210 -73 -203 -71
rect -210 -75 -208 -73
rect -206 -75 -203 -73
rect -210 -77 -203 -75
rect -201 -67 -195 -65
rect -201 -73 -193 -67
rect -201 -75 -198 -73
rect -196 -75 -193 -73
rect -201 -77 -193 -75
rect -191 -73 -183 -67
rect -191 -75 -188 -73
rect -186 -75 -183 -73
rect -191 -77 -183 -75
rect -181 -69 -174 -67
rect -181 -71 -178 -69
rect -176 -71 -174 -69
rect -165 -71 -160 -65
rect -181 -77 -174 -71
rect -167 -73 -160 -71
rect -167 -75 -165 -73
rect -163 -75 -160 -73
rect -167 -77 -160 -75
rect -158 -67 -152 -65
rect -158 -73 -150 -67
rect -158 -75 -155 -73
rect -153 -75 -150 -73
rect -158 -77 -150 -75
rect -148 -73 -140 -67
rect -148 -75 -145 -73
rect -143 -75 -140 -73
rect -148 -77 -140 -75
rect -138 -69 -131 -67
rect -138 -71 -135 -69
rect -133 -71 -131 -69
rect -122 -71 -117 -65
rect -138 -77 -131 -71
rect -124 -73 -117 -71
rect -124 -75 -122 -73
rect -120 -75 -117 -73
rect -124 -77 -117 -75
rect -115 -67 -109 -65
rect -115 -73 -107 -67
rect -115 -75 -112 -73
rect -110 -75 -107 -73
rect -115 -77 -107 -75
rect -105 -73 -97 -67
rect -105 -75 -102 -73
rect -100 -75 -97 -73
rect -105 -77 -97 -75
rect -95 -69 -88 -67
rect -95 -71 -92 -69
rect -90 -71 -88 -69
rect -95 -77 -88 -71
rect -252 -157 -247 -145
rect -254 -159 -247 -157
rect -254 -161 -252 -159
rect -250 -161 -247 -159
rect -254 -166 -247 -161
rect -254 -168 -252 -166
rect -250 -168 -247 -166
rect -254 -170 -247 -168
rect -245 -147 -236 -145
rect -245 -149 -241 -147
rect -239 -149 -236 -147
rect -213 -147 -199 -145
rect -213 -148 -206 -147
rect -245 -157 -236 -149
rect -229 -157 -224 -148
rect -245 -170 -234 -157
rect -232 -166 -224 -157
rect -232 -168 -229 -166
rect -227 -168 -224 -166
rect -232 -170 -224 -168
rect -229 -173 -224 -170
rect -222 -173 -217 -148
rect -215 -149 -206 -148
rect -204 -149 -199 -147
rect -215 -154 -199 -149
rect -215 -156 -206 -154
rect -204 -156 -199 -154
rect -215 -173 -199 -156
rect -197 -155 -189 -145
rect -197 -157 -194 -155
rect -192 -157 -189 -155
rect -197 -162 -189 -157
rect -197 -164 -194 -162
rect -192 -164 -189 -162
rect -197 -173 -189 -164
rect -187 -147 -179 -145
rect -187 -149 -184 -147
rect -182 -149 -179 -147
rect -187 -154 -179 -149
rect -187 -156 -184 -154
rect -182 -156 -179 -154
rect -187 -173 -179 -156
rect -177 -160 -172 -145
rect -150 -160 -145 -145
rect -177 -162 -170 -160
rect -177 -164 -174 -162
rect -172 -164 -170 -162
rect -177 -169 -170 -164
rect -177 -171 -174 -169
rect -172 -171 -170 -169
rect -177 -173 -170 -171
rect -152 -162 -145 -160
rect -152 -164 -150 -162
rect -148 -164 -145 -162
rect -152 -169 -145 -164
rect -152 -171 -150 -169
rect -148 -171 -145 -169
rect -152 -173 -145 -171
rect -143 -147 -135 -145
rect -143 -149 -140 -147
rect -138 -149 -135 -147
rect -143 -154 -135 -149
rect -143 -156 -140 -154
rect -138 -156 -135 -154
rect -143 -173 -135 -156
rect -133 -155 -125 -145
rect -133 -157 -130 -155
rect -128 -157 -125 -155
rect -133 -162 -125 -157
rect -133 -164 -130 -162
rect -128 -164 -125 -162
rect -133 -173 -125 -164
rect -123 -147 -109 -145
rect -123 -149 -118 -147
rect -116 -148 -109 -147
rect -86 -147 -77 -145
rect -116 -149 -107 -148
rect -123 -154 -107 -149
rect -123 -156 -118 -154
rect -116 -156 -107 -154
rect -123 -173 -107 -156
rect -105 -173 -100 -148
rect -98 -157 -93 -148
rect -86 -149 -83 -147
rect -81 -149 -77 -147
rect -86 -157 -77 -149
rect -98 -166 -90 -157
rect -98 -168 -95 -166
rect -93 -168 -90 -166
rect -98 -170 -90 -168
rect -88 -170 -77 -157
rect -75 -157 -70 -145
rect -75 -159 -68 -157
rect -75 -161 -72 -159
rect -70 -161 -68 -159
rect -75 -166 -68 -161
rect -75 -168 -72 -166
rect -70 -168 -68 -166
rect -75 -170 -68 -168
rect -98 -173 -93 -170
rect -250 -323 -245 -317
rect -252 -325 -245 -323
rect -252 -327 -250 -325
rect -248 -327 -245 -325
rect -252 -329 -245 -327
rect -243 -319 -237 -317
rect -243 -325 -235 -319
rect -243 -327 -240 -325
rect -238 -327 -235 -325
rect -243 -329 -235 -327
rect -233 -325 -225 -319
rect -233 -327 -230 -325
rect -228 -327 -225 -325
rect -233 -329 -225 -327
rect -223 -321 -216 -319
rect -223 -323 -220 -321
rect -218 -323 -216 -321
rect -207 -323 -202 -317
rect -223 -329 -216 -323
rect -209 -325 -202 -323
rect -209 -327 -207 -325
rect -205 -327 -202 -325
rect -209 -329 -202 -327
rect -200 -319 -194 -317
rect -200 -325 -192 -319
rect -200 -327 -197 -325
rect -195 -327 -192 -325
rect -200 -329 -192 -327
rect -190 -325 -182 -319
rect -190 -327 -187 -325
rect -185 -327 -182 -325
rect -190 -329 -182 -327
rect -180 -321 -173 -319
rect -180 -323 -177 -321
rect -175 -323 -173 -321
rect -164 -323 -159 -317
rect -180 -329 -173 -323
rect -166 -325 -159 -323
rect -166 -327 -164 -325
rect -162 -327 -159 -325
rect -166 -329 -159 -327
rect -157 -319 -151 -317
rect -157 -325 -149 -319
rect -157 -327 -154 -325
rect -152 -327 -149 -325
rect -157 -329 -149 -327
rect -147 -325 -139 -319
rect -147 -327 -144 -325
rect -142 -327 -139 -325
rect -147 -329 -139 -327
rect -137 -321 -130 -319
rect -137 -323 -134 -321
rect -132 -323 -130 -321
rect -121 -323 -116 -317
rect -137 -329 -130 -323
rect -123 -325 -116 -323
rect -123 -327 -121 -325
rect -119 -327 -116 -325
rect -123 -329 -116 -327
rect -114 -319 -108 -317
rect -114 -325 -106 -319
rect -114 -327 -111 -325
rect -109 -327 -106 -325
rect -114 -329 -106 -327
rect -104 -325 -96 -319
rect -104 -327 -101 -325
rect -99 -327 -96 -325
rect -104 -329 -96 -327
rect -94 -321 -87 -319
rect -94 -323 -91 -321
rect -89 -323 -87 -321
rect -94 -329 -87 -323
rect 269 171 274 177
rect 267 169 274 171
rect 267 167 269 169
rect 271 167 274 169
rect 267 165 274 167
rect 276 175 282 177
rect 276 169 284 175
rect 276 167 279 169
rect 281 167 284 169
rect 276 165 284 167
rect 286 169 294 175
rect 286 167 289 169
rect 291 167 294 169
rect 286 165 294 167
rect 296 173 303 175
rect 296 171 299 173
rect 301 171 303 173
rect 312 171 317 177
rect 296 165 303 171
rect 310 169 317 171
rect 310 167 312 169
rect 314 167 317 169
rect 310 165 317 167
rect 319 175 325 177
rect 319 169 327 175
rect 319 167 322 169
rect 324 167 327 169
rect 319 165 327 167
rect 329 169 337 175
rect 329 167 332 169
rect 334 167 337 169
rect 329 165 337 167
rect 339 173 346 175
rect 339 171 342 173
rect 344 171 346 173
rect 355 171 360 177
rect 339 165 346 171
rect 353 169 360 171
rect 353 167 355 169
rect 357 167 360 169
rect 353 165 360 167
rect 362 175 368 177
rect 362 169 370 175
rect 362 167 365 169
rect 367 167 370 169
rect 362 165 370 167
rect 372 169 380 175
rect 372 167 375 169
rect 377 167 380 169
rect 372 165 380 167
rect 382 173 389 175
rect 382 171 385 173
rect 387 171 389 173
rect 398 171 403 177
rect 382 165 389 171
rect 396 169 403 171
rect 396 167 398 169
rect 400 167 403 169
rect 396 165 403 167
rect 405 175 411 177
rect 405 169 413 175
rect 405 167 408 169
rect 410 167 413 169
rect 405 165 413 167
rect 415 169 423 175
rect 415 167 418 169
rect 420 167 423 169
rect 415 165 423 167
rect 425 173 432 175
rect 425 171 428 173
rect 430 171 432 173
rect 425 165 432 171
rect 268 85 273 97
rect 266 83 273 85
rect 266 81 268 83
rect 270 81 273 83
rect 266 76 273 81
rect 266 74 268 76
rect 270 74 273 76
rect 266 72 273 74
rect 275 95 284 97
rect 275 93 279 95
rect 281 93 284 95
rect 307 95 321 97
rect 307 94 314 95
rect 275 85 284 93
rect 291 85 296 94
rect 275 72 286 85
rect 288 76 296 85
rect 288 74 291 76
rect 293 74 296 76
rect 288 72 296 74
rect 291 69 296 72
rect 298 69 303 94
rect 305 93 314 94
rect 316 93 321 95
rect 305 88 321 93
rect 305 86 314 88
rect 316 86 321 88
rect 305 69 321 86
rect 323 87 331 97
rect 323 85 326 87
rect 328 85 331 87
rect 323 80 331 85
rect 323 78 326 80
rect 328 78 331 80
rect 323 69 331 78
rect 333 95 341 97
rect 333 93 336 95
rect 338 93 341 95
rect 333 88 341 93
rect 333 86 336 88
rect 338 86 341 88
rect 333 69 341 86
rect 343 82 348 97
rect 370 82 375 97
rect 343 80 350 82
rect 343 78 346 80
rect 348 78 350 80
rect 343 73 350 78
rect 343 71 346 73
rect 348 71 350 73
rect 343 69 350 71
rect 368 80 375 82
rect 368 78 370 80
rect 372 78 375 80
rect 368 73 375 78
rect 368 71 370 73
rect 372 71 375 73
rect 368 69 375 71
rect 377 95 385 97
rect 377 93 380 95
rect 382 93 385 95
rect 377 88 385 93
rect 377 86 380 88
rect 382 86 385 88
rect 377 69 385 86
rect 387 87 395 97
rect 387 85 390 87
rect 392 85 395 87
rect 387 80 395 85
rect 387 78 390 80
rect 392 78 395 80
rect 387 69 395 78
rect 397 95 411 97
rect 397 93 402 95
rect 404 94 411 95
rect 434 95 443 97
rect 404 93 413 94
rect 397 88 413 93
rect 397 86 402 88
rect 404 86 413 88
rect 397 69 413 86
rect 415 69 420 94
rect 422 85 427 94
rect 434 93 437 95
rect 439 93 443 95
rect 434 85 443 93
rect 422 76 430 85
rect 422 74 425 76
rect 427 74 430 76
rect 422 72 430 74
rect 432 72 443 85
rect 445 85 450 97
rect 445 83 452 85
rect 445 81 448 83
rect 450 81 452 83
rect 445 76 452 81
rect 445 74 448 76
rect 450 74 452 76
rect 445 72 452 74
rect 422 69 427 72
rect 19 -105 24 -90
rect 17 -107 24 -105
rect 17 -109 19 -107
rect 21 -109 24 -107
rect 17 -114 24 -109
rect 17 -116 19 -114
rect 21 -116 24 -114
rect 17 -118 24 -116
rect 26 -92 34 -90
rect 26 -94 29 -92
rect 31 -94 34 -92
rect 26 -99 34 -94
rect 26 -101 29 -99
rect 31 -101 34 -99
rect 26 -118 34 -101
rect 36 -100 44 -90
rect 36 -102 39 -100
rect 41 -102 44 -100
rect 36 -107 44 -102
rect 36 -109 39 -107
rect 41 -109 44 -107
rect 36 -118 44 -109
rect 46 -92 60 -90
rect 46 -94 51 -92
rect 53 -93 60 -92
rect 83 -92 92 -90
rect 53 -94 62 -93
rect 46 -99 62 -94
rect 46 -101 51 -99
rect 53 -101 62 -99
rect 46 -118 62 -101
rect 64 -118 69 -93
rect 71 -102 76 -93
rect 83 -94 86 -92
rect 88 -94 92 -92
rect 83 -102 92 -94
rect 71 -111 79 -102
rect 71 -113 74 -111
rect 76 -113 79 -111
rect 71 -115 79 -113
rect 81 -115 92 -102
rect 94 -102 99 -90
rect 107 -97 112 -90
rect 105 -99 112 -97
rect 105 -101 107 -99
rect 109 -101 112 -99
rect 94 -104 101 -102
rect 105 -103 112 -101
rect 94 -106 97 -104
rect 99 -106 101 -104
rect 94 -111 101 -106
rect 107 -108 112 -103
rect 114 -108 119 -90
rect 121 -92 130 -90
rect 121 -94 125 -92
rect 127 -94 130 -92
rect 121 -99 130 -94
rect 121 -108 132 -99
rect 94 -113 97 -111
rect 99 -113 101 -111
rect 94 -115 101 -113
rect 71 -118 76 -115
rect 124 -111 132 -108
rect 134 -101 141 -99
rect 134 -103 137 -101
rect 139 -103 141 -101
rect 134 -105 141 -103
rect 148 -105 153 -90
rect 134 -111 139 -105
rect 146 -107 153 -105
rect 146 -109 148 -107
rect 150 -109 153 -107
rect 146 -114 153 -109
rect 146 -116 148 -114
rect 150 -116 153 -114
rect 146 -118 153 -116
rect 155 -92 163 -90
rect 155 -94 158 -92
rect 160 -94 163 -92
rect 155 -99 163 -94
rect 155 -101 158 -99
rect 160 -101 163 -99
rect 155 -118 163 -101
rect 165 -100 173 -90
rect 165 -102 168 -100
rect 170 -102 173 -100
rect 165 -107 173 -102
rect 165 -109 168 -107
rect 170 -109 173 -107
rect 165 -118 173 -109
rect 175 -92 189 -90
rect 175 -94 180 -92
rect 182 -93 189 -92
rect 212 -92 221 -90
rect 182 -94 191 -93
rect 175 -99 191 -94
rect 175 -101 180 -99
rect 182 -101 191 -99
rect 175 -118 191 -101
rect 193 -118 198 -93
rect 200 -102 205 -93
rect 212 -94 215 -92
rect 217 -94 221 -92
rect 212 -102 221 -94
rect 200 -111 208 -102
rect 200 -113 203 -111
rect 205 -113 208 -111
rect 200 -115 208 -113
rect 210 -115 221 -102
rect 223 -102 228 -90
rect 238 -102 243 -90
rect 223 -104 230 -102
rect 223 -106 226 -104
rect 228 -106 230 -104
rect 223 -111 230 -106
rect 223 -113 226 -111
rect 228 -113 230 -111
rect 223 -115 230 -113
rect 236 -104 243 -102
rect 236 -106 238 -104
rect 240 -106 243 -104
rect 236 -111 243 -106
rect 236 -113 238 -111
rect 240 -113 243 -111
rect 236 -115 243 -113
rect 245 -92 254 -90
rect 245 -94 249 -92
rect 251 -94 254 -92
rect 277 -92 291 -90
rect 277 -93 284 -92
rect 245 -102 254 -94
rect 261 -102 266 -93
rect 245 -115 256 -102
rect 258 -111 266 -102
rect 258 -113 261 -111
rect 263 -113 266 -111
rect 258 -115 266 -113
rect 200 -118 205 -115
rect 261 -118 266 -115
rect 268 -118 273 -93
rect 275 -94 284 -93
rect 286 -94 291 -92
rect 275 -99 291 -94
rect 275 -101 284 -99
rect 286 -101 291 -99
rect 275 -118 291 -101
rect 293 -100 301 -90
rect 293 -102 296 -100
rect 298 -102 301 -100
rect 293 -107 301 -102
rect 293 -109 296 -107
rect 298 -109 301 -107
rect 293 -118 301 -109
rect 303 -92 311 -90
rect 303 -94 306 -92
rect 308 -94 311 -92
rect 303 -99 311 -94
rect 303 -101 306 -99
rect 308 -101 311 -99
rect 303 -118 311 -101
rect 313 -105 318 -90
rect 336 -92 345 -90
rect 336 -94 339 -92
rect 341 -94 345 -92
rect 336 -99 345 -94
rect 325 -101 332 -99
rect 325 -103 327 -101
rect 329 -103 332 -101
rect 325 -105 332 -103
rect 313 -107 320 -105
rect 313 -109 316 -107
rect 318 -109 320 -107
rect 313 -114 320 -109
rect 327 -111 332 -105
rect 334 -108 345 -99
rect 347 -108 352 -90
rect 354 -97 359 -90
rect 354 -99 361 -97
rect 354 -101 357 -99
rect 359 -101 361 -99
rect 354 -103 361 -101
rect 367 -102 372 -90
rect 354 -108 359 -103
rect 365 -104 372 -102
rect 365 -106 367 -104
rect 369 -106 372 -104
rect 334 -111 342 -108
rect 313 -116 316 -114
rect 318 -116 320 -114
rect 313 -118 320 -116
rect 365 -111 372 -106
rect 365 -113 367 -111
rect 369 -113 372 -111
rect 365 -115 372 -113
rect 374 -92 383 -90
rect 374 -94 378 -92
rect 380 -94 383 -92
rect 406 -92 420 -90
rect 406 -93 413 -92
rect 374 -102 383 -94
rect 390 -102 395 -93
rect 374 -115 385 -102
rect 387 -111 395 -102
rect 387 -113 390 -111
rect 392 -113 395 -111
rect 387 -115 395 -113
rect 390 -118 395 -115
rect 397 -118 402 -93
rect 404 -94 413 -93
rect 415 -94 420 -92
rect 404 -99 420 -94
rect 404 -101 413 -99
rect 415 -101 420 -99
rect 404 -118 420 -101
rect 422 -100 430 -90
rect 422 -102 425 -100
rect 427 -102 430 -100
rect 422 -107 430 -102
rect 422 -109 425 -107
rect 427 -109 430 -107
rect 422 -118 430 -109
rect 432 -92 440 -90
rect 432 -94 435 -92
rect 437 -94 440 -92
rect 432 -99 440 -94
rect 432 -101 435 -99
rect 437 -101 440 -99
rect 432 -118 440 -101
rect 442 -105 447 -90
rect 457 -105 462 -90
rect 442 -107 449 -105
rect 442 -109 445 -107
rect 447 -109 449 -107
rect 442 -114 449 -109
rect 442 -116 445 -114
rect 447 -116 449 -114
rect 442 -118 449 -116
rect 455 -107 462 -105
rect 455 -109 457 -107
rect 459 -109 462 -107
rect 455 -114 462 -109
rect 455 -116 457 -114
rect 459 -116 462 -114
rect 455 -118 462 -116
rect 464 -92 472 -90
rect 464 -94 467 -92
rect 469 -94 472 -92
rect 464 -99 472 -94
rect 464 -101 467 -99
rect 469 -101 472 -99
rect 464 -118 472 -101
rect 474 -100 482 -90
rect 474 -102 477 -100
rect 479 -102 482 -100
rect 474 -107 482 -102
rect 474 -109 477 -107
rect 479 -109 482 -107
rect 474 -118 482 -109
rect 484 -92 498 -90
rect 484 -94 489 -92
rect 491 -93 498 -92
rect 521 -92 530 -90
rect 491 -94 500 -93
rect 484 -99 500 -94
rect 484 -101 489 -99
rect 491 -101 500 -99
rect 484 -118 500 -101
rect 502 -118 507 -93
rect 509 -102 514 -93
rect 521 -94 524 -92
rect 526 -94 530 -92
rect 521 -102 530 -94
rect 509 -111 517 -102
rect 509 -113 512 -111
rect 514 -113 517 -111
rect 509 -115 517 -113
rect 519 -115 530 -102
rect 532 -102 537 -90
rect 545 -97 550 -90
rect 543 -99 550 -97
rect 543 -101 545 -99
rect 547 -101 550 -99
rect 532 -104 539 -102
rect 543 -103 550 -101
rect 532 -106 535 -104
rect 537 -106 539 -104
rect 532 -111 539 -106
rect 545 -108 550 -103
rect 552 -108 557 -90
rect 559 -92 568 -90
rect 559 -94 563 -92
rect 565 -94 568 -92
rect 559 -99 568 -94
rect 559 -108 570 -99
rect 532 -113 535 -111
rect 537 -113 539 -111
rect 532 -115 539 -113
rect 509 -118 514 -115
rect 562 -111 570 -108
rect 572 -101 579 -99
rect 572 -103 575 -101
rect 577 -103 579 -101
rect 572 -105 579 -103
rect 586 -105 591 -90
rect 572 -111 577 -105
rect 584 -107 591 -105
rect 584 -109 586 -107
rect 588 -109 591 -107
rect 584 -114 591 -109
rect 584 -116 586 -114
rect 588 -116 591 -114
rect 584 -118 591 -116
rect 593 -92 601 -90
rect 593 -94 596 -92
rect 598 -94 601 -92
rect 593 -99 601 -94
rect 593 -101 596 -99
rect 598 -101 601 -99
rect 593 -118 601 -101
rect 603 -100 611 -90
rect 603 -102 606 -100
rect 608 -102 611 -100
rect 603 -107 611 -102
rect 603 -109 606 -107
rect 608 -109 611 -107
rect 603 -118 611 -109
rect 613 -92 627 -90
rect 613 -94 618 -92
rect 620 -93 627 -92
rect 650 -92 659 -90
rect 620 -94 629 -93
rect 613 -99 629 -94
rect 613 -101 618 -99
rect 620 -101 629 -99
rect 613 -118 629 -101
rect 631 -118 636 -93
rect 638 -102 643 -93
rect 650 -94 653 -92
rect 655 -94 659 -92
rect 650 -102 659 -94
rect 638 -111 646 -102
rect 638 -113 641 -111
rect 643 -113 646 -111
rect 638 -115 646 -113
rect 648 -115 659 -102
rect 661 -102 666 -90
rect 661 -104 668 -102
rect 661 -106 664 -104
rect 666 -106 668 -104
rect 678 -105 683 -90
rect 661 -111 668 -106
rect 661 -113 664 -111
rect 666 -113 668 -111
rect 661 -115 668 -113
rect 676 -107 683 -105
rect 676 -109 678 -107
rect 680 -109 683 -107
rect 676 -114 683 -109
rect 638 -118 643 -115
rect 676 -116 678 -114
rect 680 -116 683 -114
rect 676 -118 683 -116
rect 685 -92 693 -90
rect 685 -94 688 -92
rect 690 -94 693 -92
rect 685 -99 693 -94
rect 685 -101 688 -99
rect 690 -101 693 -99
rect 685 -118 693 -101
rect 695 -100 703 -90
rect 695 -102 698 -100
rect 700 -102 703 -100
rect 695 -107 703 -102
rect 695 -109 698 -107
rect 700 -109 703 -107
rect 695 -118 703 -109
rect 705 -92 719 -90
rect 705 -94 710 -92
rect 712 -93 719 -92
rect 742 -92 751 -90
rect 712 -94 721 -93
rect 705 -99 721 -94
rect 705 -101 710 -99
rect 712 -101 721 -99
rect 705 -118 721 -101
rect 723 -118 728 -93
rect 730 -102 735 -93
rect 742 -94 745 -92
rect 747 -94 751 -92
rect 742 -102 751 -94
rect 730 -111 738 -102
rect 730 -113 733 -111
rect 735 -113 738 -111
rect 730 -115 738 -113
rect 740 -115 751 -102
rect 753 -102 758 -90
rect 753 -104 760 -102
rect 753 -106 756 -104
rect 758 -106 760 -104
rect 753 -111 760 -106
rect 753 -113 756 -111
rect 758 -113 760 -111
rect 753 -115 760 -113
rect 730 -118 735 -115
rect 402 -246 407 -240
rect 400 -248 407 -246
rect 400 -250 402 -248
rect 404 -250 407 -248
rect 400 -252 407 -250
rect 409 -242 415 -240
rect 409 -248 417 -242
rect 409 -250 412 -248
rect 414 -250 417 -248
rect 409 -252 417 -250
rect 419 -248 427 -242
rect 419 -250 422 -248
rect 424 -250 427 -248
rect 419 -252 427 -250
rect 429 -244 436 -242
rect 429 -246 432 -244
rect 434 -246 436 -244
rect 445 -246 450 -240
rect 429 -252 436 -246
rect 443 -248 450 -246
rect 443 -250 445 -248
rect 447 -250 450 -248
rect 443 -252 450 -250
rect 452 -242 458 -240
rect 452 -248 460 -242
rect 452 -250 455 -248
rect 457 -250 460 -248
rect 452 -252 460 -250
rect 462 -248 470 -242
rect 462 -250 465 -248
rect 467 -250 470 -248
rect 462 -252 470 -250
rect 472 -244 479 -242
rect 472 -246 475 -244
rect 477 -246 479 -244
rect 488 -246 493 -240
rect 472 -252 479 -246
rect 486 -248 493 -246
rect 486 -250 488 -248
rect 490 -250 493 -248
rect 486 -252 493 -250
rect 495 -242 501 -240
rect 495 -248 503 -242
rect 495 -250 498 -248
rect 500 -250 503 -248
rect 495 -252 503 -250
rect 505 -248 513 -242
rect 505 -250 508 -248
rect 510 -250 513 -248
rect 505 -252 513 -250
rect 515 -244 522 -242
rect 515 -246 518 -244
rect 520 -246 522 -244
rect 531 -246 536 -240
rect 515 -252 522 -246
rect 529 -248 536 -246
rect 529 -250 531 -248
rect 533 -250 536 -248
rect 529 -252 536 -250
rect 538 -242 544 -240
rect 538 -248 546 -242
rect 538 -250 541 -248
rect 543 -250 546 -248
rect 538 -252 546 -250
rect 548 -248 556 -242
rect 548 -250 551 -248
rect 553 -250 556 -248
rect 548 -252 556 -250
rect 558 -244 565 -242
rect 558 -246 561 -244
rect 563 -246 565 -244
rect 558 -252 565 -246
rect 401 -332 406 -320
rect 399 -334 406 -332
rect 399 -336 401 -334
rect 403 -336 406 -334
rect 399 -341 406 -336
rect 399 -343 401 -341
rect 403 -343 406 -341
rect 399 -345 406 -343
rect 408 -322 417 -320
rect 408 -324 412 -322
rect 414 -324 417 -322
rect 440 -322 454 -320
rect 440 -323 447 -322
rect 408 -332 417 -324
rect 424 -332 429 -323
rect 408 -345 419 -332
rect 421 -341 429 -332
rect 421 -343 424 -341
rect 426 -343 429 -341
rect 421 -345 429 -343
rect 424 -348 429 -345
rect 431 -348 436 -323
rect 438 -324 447 -323
rect 449 -324 454 -322
rect 438 -329 454 -324
rect 438 -331 447 -329
rect 449 -331 454 -329
rect 438 -348 454 -331
rect 456 -330 464 -320
rect 456 -332 459 -330
rect 461 -332 464 -330
rect 456 -337 464 -332
rect 456 -339 459 -337
rect 461 -339 464 -337
rect 456 -348 464 -339
rect 466 -322 474 -320
rect 466 -324 469 -322
rect 471 -324 474 -322
rect 466 -329 474 -324
rect 466 -331 469 -329
rect 471 -331 474 -329
rect 466 -348 474 -331
rect 476 -335 481 -320
rect 503 -335 508 -320
rect 476 -337 483 -335
rect 476 -339 479 -337
rect 481 -339 483 -337
rect 476 -344 483 -339
rect 476 -346 479 -344
rect 481 -346 483 -344
rect 476 -348 483 -346
rect 501 -337 508 -335
rect 501 -339 503 -337
rect 505 -339 508 -337
rect 501 -344 508 -339
rect 501 -346 503 -344
rect 505 -346 508 -344
rect 501 -348 508 -346
rect 510 -322 518 -320
rect 510 -324 513 -322
rect 515 -324 518 -322
rect 510 -329 518 -324
rect 510 -331 513 -329
rect 515 -331 518 -329
rect 510 -348 518 -331
rect 520 -330 528 -320
rect 520 -332 523 -330
rect 525 -332 528 -330
rect 520 -337 528 -332
rect 520 -339 523 -337
rect 525 -339 528 -337
rect 520 -348 528 -339
rect 530 -322 544 -320
rect 530 -324 535 -322
rect 537 -323 544 -322
rect 567 -322 576 -320
rect 537 -324 546 -323
rect 530 -329 546 -324
rect 530 -331 535 -329
rect 537 -331 546 -329
rect 530 -348 546 -331
rect 548 -348 553 -323
rect 555 -332 560 -323
rect 567 -324 570 -322
rect 572 -324 576 -322
rect 567 -332 576 -324
rect 555 -341 563 -332
rect 555 -343 558 -341
rect 560 -343 563 -341
rect 555 -345 563 -343
rect 565 -345 576 -332
rect 578 -332 583 -320
rect 578 -334 585 -332
rect 578 -336 581 -334
rect 583 -336 585 -334
rect 578 -341 585 -336
rect 578 -343 581 -341
rect 583 -343 585 -341
rect 578 -345 585 -343
rect 555 -348 560 -345
rect -251 -409 -246 -397
rect -253 -411 -246 -409
rect -253 -413 -251 -411
rect -249 -413 -246 -411
rect -253 -418 -246 -413
rect -253 -420 -251 -418
rect -249 -420 -246 -418
rect -253 -422 -246 -420
rect -244 -399 -235 -397
rect -244 -401 -240 -399
rect -238 -401 -235 -399
rect -212 -399 -198 -397
rect -212 -400 -205 -399
rect -244 -409 -235 -401
rect -228 -409 -223 -400
rect -244 -422 -233 -409
rect -231 -418 -223 -409
rect -231 -420 -228 -418
rect -226 -420 -223 -418
rect -231 -422 -223 -420
rect -228 -425 -223 -422
rect -221 -425 -216 -400
rect -214 -401 -205 -400
rect -203 -401 -198 -399
rect -214 -406 -198 -401
rect -214 -408 -205 -406
rect -203 -408 -198 -406
rect -214 -425 -198 -408
rect -196 -407 -188 -397
rect -196 -409 -193 -407
rect -191 -409 -188 -407
rect -196 -414 -188 -409
rect -196 -416 -193 -414
rect -191 -416 -188 -414
rect -196 -425 -188 -416
rect -186 -399 -178 -397
rect -186 -401 -183 -399
rect -181 -401 -178 -399
rect -186 -406 -178 -401
rect -186 -408 -183 -406
rect -181 -408 -178 -406
rect -186 -425 -178 -408
rect -176 -412 -171 -397
rect -149 -412 -144 -397
rect -176 -414 -169 -412
rect -176 -416 -173 -414
rect -171 -416 -169 -414
rect -176 -421 -169 -416
rect -176 -423 -173 -421
rect -171 -423 -169 -421
rect -176 -425 -169 -423
rect -151 -414 -144 -412
rect -151 -416 -149 -414
rect -147 -416 -144 -414
rect -151 -421 -144 -416
rect -151 -423 -149 -421
rect -147 -423 -144 -421
rect -151 -425 -144 -423
rect -142 -399 -134 -397
rect -142 -401 -139 -399
rect -137 -401 -134 -399
rect -142 -406 -134 -401
rect -142 -408 -139 -406
rect -137 -408 -134 -406
rect -142 -425 -134 -408
rect -132 -407 -124 -397
rect -132 -409 -129 -407
rect -127 -409 -124 -407
rect -132 -414 -124 -409
rect -132 -416 -129 -414
rect -127 -416 -124 -414
rect -132 -425 -124 -416
rect -122 -399 -108 -397
rect -122 -401 -117 -399
rect -115 -400 -108 -399
rect -85 -399 -76 -397
rect -115 -401 -106 -400
rect -122 -406 -106 -401
rect -122 -408 -117 -406
rect -115 -408 -106 -406
rect -122 -425 -106 -408
rect -104 -425 -99 -400
rect -97 -409 -92 -400
rect -85 -401 -82 -399
rect -80 -401 -76 -399
rect -85 -409 -76 -401
rect -97 -418 -89 -409
rect -97 -420 -94 -418
rect -92 -420 -89 -418
rect -97 -422 -89 -420
rect -87 -422 -76 -409
rect -74 -409 -69 -397
rect -74 -411 -67 -409
rect -74 -413 -71 -411
rect -69 -413 -67 -411
rect -74 -418 -67 -413
rect -74 -420 -71 -418
rect -69 -420 -67 -418
rect -74 -422 -67 -420
rect -97 -425 -92 -422
rect 21 -490 26 -475
rect 19 -492 26 -490
rect 19 -494 21 -492
rect 23 -494 26 -492
rect 19 -499 26 -494
rect 19 -501 21 -499
rect 23 -501 26 -499
rect 19 -503 26 -501
rect 28 -477 36 -475
rect 28 -479 31 -477
rect 33 -479 36 -477
rect 28 -484 36 -479
rect 28 -486 31 -484
rect 33 -486 36 -484
rect 28 -503 36 -486
rect 38 -485 46 -475
rect 38 -487 41 -485
rect 43 -487 46 -485
rect 38 -492 46 -487
rect 38 -494 41 -492
rect 43 -494 46 -492
rect 38 -503 46 -494
rect 48 -477 62 -475
rect 48 -479 53 -477
rect 55 -478 62 -477
rect 85 -477 94 -475
rect 55 -479 64 -478
rect 48 -484 64 -479
rect 48 -486 53 -484
rect 55 -486 64 -484
rect 48 -503 64 -486
rect 66 -503 71 -478
rect 73 -487 78 -478
rect 85 -479 88 -477
rect 90 -479 94 -477
rect 85 -487 94 -479
rect 73 -496 81 -487
rect 73 -498 76 -496
rect 78 -498 81 -496
rect 73 -500 81 -498
rect 83 -500 94 -487
rect 96 -487 101 -475
rect 109 -482 114 -475
rect 107 -484 114 -482
rect 107 -486 109 -484
rect 111 -486 114 -484
rect 96 -489 103 -487
rect 107 -488 114 -486
rect 96 -491 99 -489
rect 101 -491 103 -489
rect 96 -496 103 -491
rect 109 -493 114 -488
rect 116 -493 121 -475
rect 123 -477 132 -475
rect 123 -479 127 -477
rect 129 -479 132 -477
rect 123 -484 132 -479
rect 123 -493 134 -484
rect 96 -498 99 -496
rect 101 -498 103 -496
rect 96 -500 103 -498
rect 73 -503 78 -500
rect 126 -496 134 -493
rect 136 -486 143 -484
rect 136 -488 139 -486
rect 141 -488 143 -486
rect 136 -490 143 -488
rect 150 -490 155 -475
rect 136 -496 141 -490
rect 148 -492 155 -490
rect 148 -494 150 -492
rect 152 -494 155 -492
rect 148 -499 155 -494
rect 148 -501 150 -499
rect 152 -501 155 -499
rect 148 -503 155 -501
rect 157 -477 165 -475
rect 157 -479 160 -477
rect 162 -479 165 -477
rect 157 -484 165 -479
rect 157 -486 160 -484
rect 162 -486 165 -484
rect 157 -503 165 -486
rect 167 -485 175 -475
rect 167 -487 170 -485
rect 172 -487 175 -485
rect 167 -492 175 -487
rect 167 -494 170 -492
rect 172 -494 175 -492
rect 167 -503 175 -494
rect 177 -477 191 -475
rect 177 -479 182 -477
rect 184 -478 191 -477
rect 214 -477 223 -475
rect 184 -479 193 -478
rect 177 -484 193 -479
rect 177 -486 182 -484
rect 184 -486 193 -484
rect 177 -503 193 -486
rect 195 -503 200 -478
rect 202 -487 207 -478
rect 214 -479 217 -477
rect 219 -479 223 -477
rect 214 -487 223 -479
rect 202 -496 210 -487
rect 202 -498 205 -496
rect 207 -498 210 -496
rect 202 -500 210 -498
rect 212 -500 223 -487
rect 225 -487 230 -475
rect 240 -487 245 -475
rect 225 -489 232 -487
rect 225 -491 228 -489
rect 230 -491 232 -489
rect 225 -496 232 -491
rect 225 -498 228 -496
rect 230 -498 232 -496
rect 225 -500 232 -498
rect 238 -489 245 -487
rect 238 -491 240 -489
rect 242 -491 245 -489
rect 238 -496 245 -491
rect 238 -498 240 -496
rect 242 -498 245 -496
rect 238 -500 245 -498
rect 247 -477 256 -475
rect 247 -479 251 -477
rect 253 -479 256 -477
rect 279 -477 293 -475
rect 279 -478 286 -477
rect 247 -487 256 -479
rect 263 -487 268 -478
rect 247 -500 258 -487
rect 260 -496 268 -487
rect 260 -498 263 -496
rect 265 -498 268 -496
rect 260 -500 268 -498
rect 202 -503 207 -500
rect 263 -503 268 -500
rect 270 -503 275 -478
rect 277 -479 286 -478
rect 288 -479 293 -477
rect 277 -484 293 -479
rect 277 -486 286 -484
rect 288 -486 293 -484
rect 277 -503 293 -486
rect 295 -485 303 -475
rect 295 -487 298 -485
rect 300 -487 303 -485
rect 295 -492 303 -487
rect 295 -494 298 -492
rect 300 -494 303 -492
rect 295 -503 303 -494
rect 305 -477 313 -475
rect 305 -479 308 -477
rect 310 -479 313 -477
rect 305 -484 313 -479
rect 305 -486 308 -484
rect 310 -486 313 -484
rect 305 -503 313 -486
rect 315 -490 320 -475
rect 338 -477 347 -475
rect 338 -479 341 -477
rect 343 -479 347 -477
rect 338 -484 347 -479
rect 327 -486 334 -484
rect 327 -488 329 -486
rect 331 -488 334 -486
rect 327 -490 334 -488
rect 315 -492 322 -490
rect 315 -494 318 -492
rect 320 -494 322 -492
rect 315 -499 322 -494
rect 329 -496 334 -490
rect 336 -493 347 -484
rect 349 -493 354 -475
rect 356 -482 361 -475
rect 356 -484 363 -482
rect 356 -486 359 -484
rect 361 -486 363 -484
rect 356 -488 363 -486
rect 369 -487 374 -475
rect 356 -493 361 -488
rect 367 -489 374 -487
rect 367 -491 369 -489
rect 371 -491 374 -489
rect 336 -496 344 -493
rect 315 -501 318 -499
rect 320 -501 322 -499
rect 315 -503 322 -501
rect 367 -496 374 -491
rect 367 -498 369 -496
rect 371 -498 374 -496
rect 367 -500 374 -498
rect 376 -477 385 -475
rect 376 -479 380 -477
rect 382 -479 385 -477
rect 408 -477 422 -475
rect 408 -478 415 -477
rect 376 -487 385 -479
rect 392 -487 397 -478
rect 376 -500 387 -487
rect 389 -496 397 -487
rect 389 -498 392 -496
rect 394 -498 397 -496
rect 389 -500 397 -498
rect 392 -503 397 -500
rect 399 -503 404 -478
rect 406 -479 415 -478
rect 417 -479 422 -477
rect 406 -484 422 -479
rect 406 -486 415 -484
rect 417 -486 422 -484
rect 406 -503 422 -486
rect 424 -485 432 -475
rect 424 -487 427 -485
rect 429 -487 432 -485
rect 424 -492 432 -487
rect 424 -494 427 -492
rect 429 -494 432 -492
rect 424 -503 432 -494
rect 434 -477 442 -475
rect 434 -479 437 -477
rect 439 -479 442 -477
rect 434 -484 442 -479
rect 434 -486 437 -484
rect 439 -486 442 -484
rect 434 -503 442 -486
rect 444 -490 449 -475
rect 459 -490 464 -475
rect 444 -492 451 -490
rect 444 -494 447 -492
rect 449 -494 451 -492
rect 444 -499 451 -494
rect 444 -501 447 -499
rect 449 -501 451 -499
rect 444 -503 451 -501
rect 457 -492 464 -490
rect 457 -494 459 -492
rect 461 -494 464 -492
rect 457 -499 464 -494
rect 457 -501 459 -499
rect 461 -501 464 -499
rect 457 -503 464 -501
rect 466 -477 474 -475
rect 466 -479 469 -477
rect 471 -479 474 -477
rect 466 -484 474 -479
rect 466 -486 469 -484
rect 471 -486 474 -484
rect 466 -503 474 -486
rect 476 -485 484 -475
rect 476 -487 479 -485
rect 481 -487 484 -485
rect 476 -492 484 -487
rect 476 -494 479 -492
rect 481 -494 484 -492
rect 476 -503 484 -494
rect 486 -477 500 -475
rect 486 -479 491 -477
rect 493 -478 500 -477
rect 523 -477 532 -475
rect 493 -479 502 -478
rect 486 -484 502 -479
rect 486 -486 491 -484
rect 493 -486 502 -484
rect 486 -503 502 -486
rect 504 -503 509 -478
rect 511 -487 516 -478
rect 523 -479 526 -477
rect 528 -479 532 -477
rect 523 -487 532 -479
rect 511 -496 519 -487
rect 511 -498 514 -496
rect 516 -498 519 -496
rect 511 -500 519 -498
rect 521 -500 532 -487
rect 534 -487 539 -475
rect 547 -482 552 -475
rect 545 -484 552 -482
rect 545 -486 547 -484
rect 549 -486 552 -484
rect 534 -489 541 -487
rect 545 -488 552 -486
rect 534 -491 537 -489
rect 539 -491 541 -489
rect 534 -496 541 -491
rect 547 -493 552 -488
rect 554 -493 559 -475
rect 561 -477 570 -475
rect 561 -479 565 -477
rect 567 -479 570 -477
rect 561 -484 570 -479
rect 561 -493 572 -484
rect 534 -498 537 -496
rect 539 -498 541 -496
rect 534 -500 541 -498
rect 511 -503 516 -500
rect 564 -496 572 -493
rect 574 -486 581 -484
rect 574 -488 577 -486
rect 579 -488 581 -486
rect 574 -490 581 -488
rect 588 -490 593 -475
rect 574 -496 579 -490
rect 586 -492 593 -490
rect 586 -494 588 -492
rect 590 -494 593 -492
rect 586 -499 593 -494
rect 586 -501 588 -499
rect 590 -501 593 -499
rect 586 -503 593 -501
rect 595 -477 603 -475
rect 595 -479 598 -477
rect 600 -479 603 -477
rect 595 -484 603 -479
rect 595 -486 598 -484
rect 600 -486 603 -484
rect 595 -503 603 -486
rect 605 -485 613 -475
rect 605 -487 608 -485
rect 610 -487 613 -485
rect 605 -492 613 -487
rect 605 -494 608 -492
rect 610 -494 613 -492
rect 605 -503 613 -494
rect 615 -477 629 -475
rect 615 -479 620 -477
rect 622 -478 629 -477
rect 652 -477 661 -475
rect 622 -479 631 -478
rect 615 -484 631 -479
rect 615 -486 620 -484
rect 622 -486 631 -484
rect 615 -503 631 -486
rect 633 -503 638 -478
rect 640 -487 645 -478
rect 652 -479 655 -477
rect 657 -479 661 -477
rect 652 -487 661 -479
rect 640 -496 648 -487
rect 640 -498 643 -496
rect 645 -498 648 -496
rect 640 -500 648 -498
rect 650 -500 661 -487
rect 663 -487 668 -475
rect 663 -489 670 -487
rect 663 -491 666 -489
rect 668 -491 670 -489
rect 680 -490 685 -475
rect 663 -496 670 -491
rect 663 -498 666 -496
rect 668 -498 670 -496
rect 663 -500 670 -498
rect 678 -492 685 -490
rect 678 -494 680 -492
rect 682 -494 685 -492
rect 678 -499 685 -494
rect 640 -503 645 -500
rect 678 -501 680 -499
rect 682 -501 685 -499
rect 678 -503 685 -501
rect 687 -477 695 -475
rect 687 -479 690 -477
rect 692 -479 695 -477
rect 687 -484 695 -479
rect 687 -486 690 -484
rect 692 -486 695 -484
rect 687 -503 695 -486
rect 697 -485 705 -475
rect 697 -487 700 -485
rect 702 -487 705 -485
rect 697 -492 705 -487
rect 697 -494 700 -492
rect 702 -494 705 -492
rect 697 -503 705 -494
rect 707 -477 721 -475
rect 707 -479 712 -477
rect 714 -478 721 -477
rect 744 -477 753 -475
rect 714 -479 723 -478
rect 707 -484 723 -479
rect 707 -486 712 -484
rect 714 -486 723 -484
rect 707 -503 723 -486
rect 725 -503 730 -478
rect 732 -487 737 -478
rect 744 -479 747 -477
rect 749 -479 753 -477
rect 744 -487 753 -479
rect 732 -496 740 -487
rect 732 -498 735 -496
rect 737 -498 740 -496
rect 732 -500 740 -498
rect 742 -500 753 -487
rect 755 -487 760 -475
rect 755 -489 762 -487
rect 755 -491 758 -489
rect 760 -491 762 -489
rect 755 -496 762 -491
rect 755 -498 758 -496
rect 760 -498 762 -496
rect 755 -500 762 -498
rect 732 -503 737 -500
rect -246 -624 -241 -609
rect -248 -626 -241 -624
rect -248 -628 -246 -626
rect -244 -628 -241 -626
rect -248 -633 -241 -628
rect -248 -635 -246 -633
rect -244 -635 -241 -633
rect -248 -637 -241 -635
rect -239 -611 -231 -609
rect -239 -613 -236 -611
rect -234 -613 -231 -611
rect -239 -618 -231 -613
rect -239 -620 -236 -618
rect -234 -620 -231 -618
rect -239 -637 -231 -620
rect -229 -619 -221 -609
rect -229 -621 -226 -619
rect -224 -621 -221 -619
rect -229 -626 -221 -621
rect -229 -628 -226 -626
rect -224 -628 -221 -626
rect -229 -637 -221 -628
rect -219 -611 -205 -609
rect -219 -613 -214 -611
rect -212 -612 -205 -611
rect -182 -611 -173 -609
rect -212 -613 -203 -612
rect -219 -618 -203 -613
rect -219 -620 -214 -618
rect -212 -620 -203 -618
rect -219 -637 -203 -620
rect -201 -637 -196 -612
rect -194 -621 -189 -612
rect -182 -613 -179 -611
rect -177 -613 -173 -611
rect -182 -621 -173 -613
rect -194 -630 -186 -621
rect -194 -632 -191 -630
rect -189 -632 -186 -630
rect -194 -634 -186 -632
rect -184 -634 -173 -621
rect -171 -621 -166 -609
rect -158 -616 -153 -609
rect -160 -618 -153 -616
rect -160 -620 -158 -618
rect -156 -620 -153 -618
rect -171 -623 -164 -621
rect -160 -622 -153 -620
rect -171 -625 -168 -623
rect -166 -625 -164 -623
rect -171 -630 -164 -625
rect -158 -627 -153 -622
rect -151 -627 -146 -609
rect -144 -611 -135 -609
rect -144 -613 -140 -611
rect -138 -613 -135 -611
rect -144 -618 -135 -613
rect -144 -627 -133 -618
rect -171 -632 -168 -630
rect -166 -632 -164 -630
rect -171 -634 -164 -632
rect -194 -637 -189 -634
rect -141 -630 -133 -627
rect -131 -620 -124 -618
rect -131 -622 -128 -620
rect -126 -622 -124 -620
rect -131 -624 -124 -622
rect -117 -624 -112 -609
rect -131 -630 -126 -624
rect -119 -626 -112 -624
rect -119 -628 -117 -626
rect -115 -628 -112 -626
rect -119 -633 -112 -628
rect -119 -635 -117 -633
rect -115 -635 -112 -633
rect -119 -637 -112 -635
rect -110 -611 -102 -609
rect -110 -613 -107 -611
rect -105 -613 -102 -611
rect -110 -618 -102 -613
rect -110 -620 -107 -618
rect -105 -620 -102 -618
rect -110 -637 -102 -620
rect -100 -619 -92 -609
rect -100 -621 -97 -619
rect -95 -621 -92 -619
rect -100 -626 -92 -621
rect -100 -628 -97 -626
rect -95 -628 -92 -626
rect -100 -637 -92 -628
rect -90 -611 -76 -609
rect -90 -613 -85 -611
rect -83 -612 -76 -611
rect -53 -611 -44 -609
rect -83 -613 -74 -612
rect -90 -618 -74 -613
rect -90 -620 -85 -618
rect -83 -620 -74 -618
rect -90 -637 -74 -620
rect -72 -637 -67 -612
rect -65 -621 -60 -612
rect -53 -613 -50 -611
rect -48 -613 -44 -611
rect -53 -621 -44 -613
rect -65 -630 -57 -621
rect -65 -632 -62 -630
rect -60 -632 -57 -630
rect -65 -634 -57 -632
rect -55 -634 -44 -621
rect -42 -621 -37 -609
rect -27 -621 -22 -609
rect -42 -623 -35 -621
rect -42 -625 -39 -623
rect -37 -625 -35 -623
rect -42 -630 -35 -625
rect -42 -632 -39 -630
rect -37 -632 -35 -630
rect -42 -634 -35 -632
rect -29 -623 -22 -621
rect -29 -625 -27 -623
rect -25 -625 -22 -623
rect -29 -630 -22 -625
rect -29 -632 -27 -630
rect -25 -632 -22 -630
rect -29 -634 -22 -632
rect -20 -611 -11 -609
rect -20 -613 -16 -611
rect -14 -613 -11 -611
rect 12 -611 26 -609
rect 12 -612 19 -611
rect -20 -621 -11 -613
rect -4 -621 1 -612
rect -20 -634 -9 -621
rect -7 -630 1 -621
rect -7 -632 -4 -630
rect -2 -632 1 -630
rect -7 -634 1 -632
rect -65 -637 -60 -634
rect -4 -637 1 -634
rect 3 -637 8 -612
rect 10 -613 19 -612
rect 21 -613 26 -611
rect 10 -618 26 -613
rect 10 -620 19 -618
rect 21 -620 26 -618
rect 10 -637 26 -620
rect 28 -619 36 -609
rect 28 -621 31 -619
rect 33 -621 36 -619
rect 28 -626 36 -621
rect 28 -628 31 -626
rect 33 -628 36 -626
rect 28 -637 36 -628
rect 38 -611 46 -609
rect 38 -613 41 -611
rect 43 -613 46 -611
rect 38 -618 46 -613
rect 38 -620 41 -618
rect 43 -620 46 -618
rect 38 -637 46 -620
rect 48 -624 53 -609
rect 71 -611 80 -609
rect 71 -613 74 -611
rect 76 -613 80 -611
rect 71 -618 80 -613
rect 60 -620 67 -618
rect 60 -622 62 -620
rect 64 -622 67 -620
rect 60 -624 67 -622
rect 48 -626 55 -624
rect 48 -628 51 -626
rect 53 -628 55 -626
rect 48 -633 55 -628
rect 62 -630 67 -624
rect 69 -627 80 -618
rect 82 -627 87 -609
rect 89 -616 94 -609
rect 89 -618 96 -616
rect 89 -620 92 -618
rect 94 -620 96 -618
rect 89 -622 96 -620
rect 102 -621 107 -609
rect 89 -627 94 -622
rect 100 -623 107 -621
rect 100 -625 102 -623
rect 104 -625 107 -623
rect 69 -630 77 -627
rect 48 -635 51 -633
rect 53 -635 55 -633
rect 48 -637 55 -635
rect 100 -630 107 -625
rect 100 -632 102 -630
rect 104 -632 107 -630
rect 100 -634 107 -632
rect 109 -611 118 -609
rect 109 -613 113 -611
rect 115 -613 118 -611
rect 141 -611 155 -609
rect 141 -612 148 -611
rect 109 -621 118 -613
rect 125 -621 130 -612
rect 109 -634 120 -621
rect 122 -630 130 -621
rect 122 -632 125 -630
rect 127 -632 130 -630
rect 122 -634 130 -632
rect 125 -637 130 -634
rect 132 -637 137 -612
rect 139 -613 148 -612
rect 150 -613 155 -611
rect 139 -618 155 -613
rect 139 -620 148 -618
rect 150 -620 155 -618
rect 139 -637 155 -620
rect 157 -619 165 -609
rect 157 -621 160 -619
rect 162 -621 165 -619
rect 157 -626 165 -621
rect 157 -628 160 -626
rect 162 -628 165 -626
rect 157 -637 165 -628
rect 167 -611 175 -609
rect 167 -613 170 -611
rect 172 -613 175 -611
rect 167 -618 175 -613
rect 167 -620 170 -618
rect 172 -620 175 -618
rect 167 -637 175 -620
rect 177 -624 182 -609
rect 192 -624 197 -609
rect 177 -626 184 -624
rect 177 -628 180 -626
rect 182 -628 184 -626
rect 177 -633 184 -628
rect 177 -635 180 -633
rect 182 -635 184 -633
rect 177 -637 184 -635
rect 190 -626 197 -624
rect 190 -628 192 -626
rect 194 -628 197 -626
rect 190 -633 197 -628
rect 190 -635 192 -633
rect 194 -635 197 -633
rect 190 -637 197 -635
rect 199 -611 207 -609
rect 199 -613 202 -611
rect 204 -613 207 -611
rect 199 -618 207 -613
rect 199 -620 202 -618
rect 204 -620 207 -618
rect 199 -637 207 -620
rect 209 -619 217 -609
rect 209 -621 212 -619
rect 214 -621 217 -619
rect 209 -626 217 -621
rect 209 -628 212 -626
rect 214 -628 217 -626
rect 209 -637 217 -628
rect 219 -611 233 -609
rect 219 -613 224 -611
rect 226 -612 233 -611
rect 256 -611 265 -609
rect 226 -613 235 -612
rect 219 -618 235 -613
rect 219 -620 224 -618
rect 226 -620 235 -618
rect 219 -637 235 -620
rect 237 -637 242 -612
rect 244 -621 249 -612
rect 256 -613 259 -611
rect 261 -613 265 -611
rect 256 -621 265 -613
rect 244 -630 252 -621
rect 244 -632 247 -630
rect 249 -632 252 -630
rect 244 -634 252 -632
rect 254 -634 265 -621
rect 267 -621 272 -609
rect 280 -616 285 -609
rect 278 -618 285 -616
rect 278 -620 280 -618
rect 282 -620 285 -618
rect 267 -623 274 -621
rect 278 -622 285 -620
rect 267 -625 270 -623
rect 272 -625 274 -623
rect 267 -630 274 -625
rect 280 -627 285 -622
rect 287 -627 292 -609
rect 294 -611 303 -609
rect 294 -613 298 -611
rect 300 -613 303 -611
rect 294 -618 303 -613
rect 294 -627 305 -618
rect 267 -632 270 -630
rect 272 -632 274 -630
rect 267 -634 274 -632
rect 244 -637 249 -634
rect 297 -630 305 -627
rect 307 -620 314 -618
rect 307 -622 310 -620
rect 312 -622 314 -620
rect 307 -624 314 -622
rect 321 -624 326 -609
rect 307 -630 312 -624
rect 319 -626 326 -624
rect 319 -628 321 -626
rect 323 -628 326 -626
rect 319 -633 326 -628
rect 319 -635 321 -633
rect 323 -635 326 -633
rect 319 -637 326 -635
rect 328 -611 336 -609
rect 328 -613 331 -611
rect 333 -613 336 -611
rect 328 -618 336 -613
rect 328 -620 331 -618
rect 333 -620 336 -618
rect 328 -637 336 -620
rect 338 -619 346 -609
rect 338 -621 341 -619
rect 343 -621 346 -619
rect 338 -626 346 -621
rect 338 -628 341 -626
rect 343 -628 346 -626
rect 338 -637 346 -628
rect 348 -611 362 -609
rect 348 -613 353 -611
rect 355 -612 362 -611
rect 385 -611 394 -609
rect 355 -613 364 -612
rect 348 -618 364 -613
rect 348 -620 353 -618
rect 355 -620 364 -618
rect 348 -637 364 -620
rect 366 -637 371 -612
rect 373 -621 378 -612
rect 385 -613 388 -611
rect 390 -613 394 -611
rect 385 -621 394 -613
rect 373 -630 381 -621
rect 373 -632 376 -630
rect 378 -632 381 -630
rect 373 -634 381 -632
rect 383 -634 394 -621
rect 396 -621 401 -609
rect 396 -623 403 -621
rect 396 -625 399 -623
rect 401 -625 403 -623
rect 413 -624 418 -609
rect 396 -630 403 -625
rect 396 -632 399 -630
rect 401 -632 403 -630
rect 396 -634 403 -632
rect 411 -626 418 -624
rect 411 -628 413 -626
rect 415 -628 418 -626
rect 411 -633 418 -628
rect 373 -637 378 -634
rect 411 -635 413 -633
rect 415 -635 418 -633
rect 411 -637 418 -635
rect 420 -611 428 -609
rect 420 -613 423 -611
rect 425 -613 428 -611
rect 420 -618 428 -613
rect 420 -620 423 -618
rect 425 -620 428 -618
rect 420 -637 428 -620
rect 430 -619 438 -609
rect 430 -621 433 -619
rect 435 -621 438 -619
rect 430 -626 438 -621
rect 430 -628 433 -626
rect 435 -628 438 -626
rect 430 -637 438 -628
rect 440 -611 454 -609
rect 440 -613 445 -611
rect 447 -612 454 -611
rect 477 -611 486 -609
rect 447 -613 456 -612
rect 440 -618 456 -613
rect 440 -620 445 -618
rect 447 -620 456 -618
rect 440 -637 456 -620
rect 458 -637 463 -612
rect 465 -621 470 -612
rect 477 -613 480 -611
rect 482 -613 486 -611
rect 477 -621 486 -613
rect 465 -630 473 -621
rect 465 -632 468 -630
rect 470 -632 473 -630
rect 465 -634 473 -632
rect 475 -634 486 -621
rect 488 -621 493 -609
rect 488 -623 495 -621
rect 488 -625 491 -623
rect 493 -625 495 -623
rect 488 -630 495 -625
rect 488 -632 491 -630
rect 493 -632 495 -630
rect 488 -634 495 -632
rect 465 -637 470 -634
<< alu1 >>
rect -336 239 874 281
rect -215 -43 -208 -38
rect -49 -43 -42 239
rect 327 199 333 239
rect 263 194 457 199
rect 263 192 270 194
rect 272 192 284 194
rect 286 192 298 194
rect 300 192 313 194
rect 315 192 327 194
rect 329 192 341 194
rect 343 192 356 194
rect 358 192 370 194
rect 372 192 384 194
rect 386 192 399 194
rect 401 192 413 194
rect 415 192 427 194
rect 429 192 457 194
rect 263 191 457 192
rect 267 169 271 178
rect 267 167 269 169
rect 267 153 271 167
rect 282 184 295 186
rect 282 182 286 184
rect 288 182 295 184
rect 282 180 295 182
rect 282 173 288 180
rect 310 169 314 178
rect 310 167 312 169
rect 267 151 268 153
rect 270 151 271 153
rect 267 146 271 151
rect 267 144 269 146
rect 271 144 279 146
rect 267 140 279 144
rect 299 153 303 162
rect 290 152 303 153
rect 290 150 295 152
rect 297 150 303 152
rect 290 148 303 150
rect 310 152 314 167
rect 325 184 333 186
rect 325 182 329 184
rect 331 182 333 184
rect 325 180 333 182
rect 325 173 331 180
rect 353 169 357 178
rect 353 167 355 169
rect 310 150 311 152
rect 313 150 314 152
rect 310 146 314 150
rect 310 144 312 146
rect 314 144 322 146
rect 310 140 322 144
rect 342 153 346 162
rect 333 152 346 153
rect 333 150 338 152
rect 340 150 346 152
rect 333 148 346 150
rect 353 152 357 167
rect 368 173 374 178
rect 396 169 400 178
rect 396 167 398 169
rect 353 150 354 152
rect 356 150 357 152
rect 353 146 357 150
rect 353 144 355 146
rect 357 144 365 146
rect 353 140 365 144
rect 385 153 389 162
rect 376 152 389 153
rect 376 150 381 152
rect 383 150 389 152
rect 376 148 389 150
rect 396 146 400 167
rect 411 184 424 186
rect 411 182 415 184
rect 417 182 424 184
rect 411 180 424 182
rect 411 173 417 180
rect 396 144 398 146
rect 400 144 408 146
rect 396 143 408 144
rect 396 141 398 143
rect 400 141 408 143
rect 396 140 408 141
rect 428 153 432 162
rect 419 152 432 153
rect 419 150 424 152
rect 426 150 432 152
rect 419 148 432 150
rect 247 134 436 135
rect 247 132 270 134
rect 272 132 280 134
rect 282 132 313 134
rect 315 132 323 134
rect 325 132 356 134
rect 358 132 366 134
rect 368 132 399 134
rect 401 132 409 134
rect 411 132 436 134
rect 247 127 436 132
rect 247 39 254 127
rect 450 103 457 191
rect 262 95 457 103
rect 266 85 279 89
rect 439 85 452 89
rect 266 83 271 85
rect 266 81 268 83
rect 270 81 271 83
rect 266 76 271 81
rect 266 74 268 76
rect 270 74 271 76
rect 266 72 271 74
rect 266 54 270 72
rect 297 72 335 73
rect 297 70 307 72
rect 309 70 335 72
rect 297 69 335 70
rect 297 66 302 69
rect 294 64 302 66
rect 294 62 295 64
rect 297 62 302 64
rect 294 60 302 62
rect 312 64 327 65
rect 312 62 314 64
rect 316 62 321 64
rect 323 62 327 64
rect 312 61 327 62
rect 314 60 318 61
rect 345 80 351 82
rect 345 78 346 80
rect 348 78 351 80
rect 345 73 351 78
rect 345 71 346 73
rect 348 71 351 73
rect 345 69 351 71
rect 314 58 315 60
rect 317 58 318 60
rect 266 52 267 54
rect 269 52 270 54
rect 266 50 270 52
rect 266 48 271 50
rect 314 52 318 58
rect 347 53 351 69
rect 367 80 373 82
rect 447 83 452 85
rect 447 81 448 83
rect 450 81 452 83
rect 367 78 370 80
rect 372 78 373 80
rect 367 73 373 78
rect 367 71 370 73
rect 372 71 373 73
rect 367 69 373 71
rect 367 61 371 69
rect 383 72 421 73
rect 383 70 417 72
rect 419 70 421 72
rect 383 69 421 70
rect 367 59 368 61
rect 370 59 371 61
rect 416 66 421 69
rect 391 64 406 65
rect 391 62 395 64
rect 397 62 402 64
rect 404 62 406 64
rect 391 61 406 62
rect 416 64 424 66
rect 416 62 421 64
rect 423 62 424 64
rect 347 52 355 53
rect 347 50 352 52
rect 354 50 355 52
rect 347 49 355 50
rect 367 49 371 59
rect 400 52 404 61
rect 416 60 424 62
rect 447 76 452 81
rect 447 74 448 76
rect 450 74 452 76
rect 447 72 452 74
rect 266 46 268 48
rect 270 46 271 48
rect 266 44 271 46
rect 329 48 351 49
rect 329 46 346 48
rect 348 46 351 48
rect 329 45 351 46
rect 367 48 389 49
rect 367 46 370 48
rect 372 46 389 48
rect 367 45 389 46
rect 448 55 452 72
rect 448 53 449 55
rect 451 53 452 55
rect 448 50 452 53
rect 447 48 452 50
rect 447 46 448 48
rect 450 46 452 48
rect 447 44 452 46
rect 247 31 790 39
rect -257 -48 -42 -43
rect -257 -50 -250 -48
rect -248 -50 -236 -48
rect -234 -50 -222 -48
rect -220 -50 -207 -48
rect -205 -50 -193 -48
rect -191 -50 -179 -48
rect -177 -50 -164 -48
rect -162 -50 -150 -48
rect -148 -50 -136 -48
rect -134 -50 -121 -48
rect -119 -50 -107 -48
rect -105 -50 -93 -48
rect -91 -50 -42 -48
rect -257 -51 -42 -50
rect -253 -73 -249 -64
rect -253 -75 -251 -73
rect -253 -89 -249 -75
rect -238 -58 -225 -56
rect -238 -60 -234 -58
rect -232 -60 -228 -58
rect -226 -60 -225 -58
rect -238 -62 -225 -60
rect -238 -69 -232 -62
rect -210 -73 -206 -64
rect -210 -75 -208 -73
rect -253 -91 -252 -89
rect -250 -91 -249 -89
rect -253 -96 -249 -91
rect -253 -98 -251 -96
rect -249 -98 -241 -96
rect -253 -102 -241 -98
rect -221 -89 -217 -80
rect -230 -90 -217 -89
rect -230 -92 -225 -90
rect -223 -92 -217 -90
rect -230 -94 -217 -92
rect -210 -90 -206 -75
rect -195 -58 -187 -56
rect -195 -60 -191 -58
rect -189 -60 -187 -58
rect -195 -62 -187 -60
rect -195 -69 -189 -62
rect -167 -73 -163 -64
rect -167 -75 -165 -73
rect -210 -92 -209 -90
rect -207 -92 -206 -90
rect -210 -96 -206 -92
rect -210 -98 -208 -96
rect -206 -98 -198 -96
rect -210 -102 -198 -98
rect -178 -89 -174 -80
rect -187 -90 -174 -89
rect -187 -92 -182 -90
rect -180 -92 -174 -90
rect -187 -94 -174 -92
rect -167 -90 -163 -75
rect -152 -69 -146 -64
rect -124 -66 -120 -64
rect -124 -68 -123 -66
rect -121 -68 -120 -66
rect -124 -73 -120 -68
rect -124 -75 -122 -73
rect -167 -92 -166 -90
rect -164 -92 -163 -90
rect -167 -96 -163 -92
rect -167 -98 -165 -96
rect -163 -98 -155 -96
rect -167 -102 -155 -98
rect -135 -89 -131 -80
rect -144 -90 -131 -89
rect -144 -92 -139 -90
rect -137 -92 -131 -90
rect -144 -94 -131 -92
rect -124 -96 -120 -75
rect -109 -57 -96 -56
rect -109 -58 -99 -57
rect -109 -60 -105 -58
rect -103 -59 -99 -58
rect -97 -59 -96 -57
rect -103 -60 -96 -59
rect -109 -62 -96 -60
rect -109 -69 -103 -62
rect -124 -98 -122 -96
rect -120 -98 -112 -96
rect -124 -102 -112 -98
rect -92 -89 -88 -80
rect -101 -90 -88 -89
rect -101 -92 -96 -90
rect -94 -92 -88 -90
rect -101 -94 -88 -92
rect -49 -84 -42 -51
rect -49 -89 765 -84
rect -49 -91 136 -89
rect 138 -91 328 -89
rect 330 -91 574 -89
rect 576 -91 765 -89
rect -284 -108 -84 -107
rect -284 -110 -250 -108
rect -248 -110 -240 -108
rect -238 -110 -207 -108
rect -205 -110 -197 -108
rect -195 -110 -164 -108
rect -162 -110 -154 -108
rect -152 -110 -121 -108
rect -119 -110 -111 -108
rect -109 -110 -84 -108
rect -284 -114 -84 -110
rect -284 -204 -278 -114
rect -257 -115 -84 -114
rect -49 -139 -42 -91
rect 14 -92 765 -91
rect 88 -102 101 -98
rect 128 -99 141 -98
rect 128 -101 129 -99
rect 131 -101 141 -99
rect 128 -102 137 -101
rect -258 -147 -42 -139
rect 16 -107 22 -105
rect 96 -104 101 -102
rect 96 -106 97 -104
rect 99 -106 101 -104
rect 16 -109 19 -107
rect 21 -109 22 -107
rect 16 -114 22 -109
rect 16 -116 19 -114
rect 21 -116 22 -114
rect 16 -118 22 -116
rect 16 -138 20 -118
rect 32 -118 70 -114
rect 65 -121 70 -118
rect 40 -123 55 -122
rect 40 -125 44 -123
rect 46 -125 51 -123
rect 53 -125 55 -123
rect 40 -126 55 -125
rect 65 -123 73 -121
rect 65 -125 66 -123
rect 68 -125 70 -123
rect 72 -125 73 -123
rect 49 -132 53 -126
rect 65 -127 73 -125
rect 96 -111 101 -106
rect 96 -113 97 -111
rect 99 -113 101 -111
rect 96 -115 101 -113
rect 97 -123 101 -115
rect 97 -125 98 -123
rect 100 -125 101 -123
rect 49 -134 50 -132
rect 52 -134 53 -132
rect 49 -135 53 -134
rect 16 -139 38 -138
rect 16 -141 19 -139
rect 21 -141 38 -139
rect 16 -142 38 -141
rect 97 -137 101 -125
rect 105 -114 109 -113
rect 105 -116 106 -114
rect 108 -116 109 -114
rect 105 -122 109 -116
rect 113 -114 117 -105
rect 139 -103 141 -101
rect 217 -102 230 -98
rect 113 -115 126 -114
rect 113 -117 120 -115
rect 122 -117 123 -115
rect 125 -117 126 -115
rect 113 -118 126 -117
rect 105 -123 118 -122
rect 105 -125 110 -123
rect 112 -125 118 -123
rect 105 -126 118 -125
rect 105 -127 109 -126
rect 96 -139 101 -137
rect 96 -141 97 -139
rect 99 -141 101 -139
rect 96 -143 101 -141
rect -254 -157 -241 -153
rect -81 -157 -68 -153
rect -254 -159 -249 -157
rect -254 -161 -252 -159
rect -250 -161 -249 -159
rect -254 -166 -249 -161
rect -254 -168 -252 -166
rect -250 -168 -249 -166
rect -254 -170 -249 -168
rect -254 -180 -250 -170
rect -223 -170 -185 -169
rect -223 -172 -213 -170
rect -211 -172 -185 -170
rect -223 -173 -185 -172
rect -254 -182 -253 -180
rect -251 -182 -250 -180
rect -254 -192 -250 -182
rect -223 -176 -218 -173
rect -226 -178 -218 -176
rect -226 -180 -225 -178
rect -223 -180 -218 -178
rect -226 -182 -218 -180
rect -208 -178 -193 -177
rect -208 -180 -206 -178
rect -204 -180 -199 -178
rect -197 -180 -193 -178
rect -208 -181 -193 -180
rect -206 -182 -202 -181
rect -175 -162 -169 -160
rect -175 -164 -174 -162
rect -172 -164 -169 -162
rect -175 -169 -169 -164
rect -175 -171 -174 -169
rect -172 -171 -169 -169
rect -175 -173 -169 -171
rect -206 -184 -205 -182
rect -203 -184 -202 -182
rect -254 -194 -249 -192
rect -206 -190 -202 -184
rect -173 -192 -169 -173
rect -153 -162 -147 -160
rect -73 -159 -68 -157
rect -73 -161 -72 -159
rect -70 -161 -68 -159
rect -153 -164 -150 -162
rect -148 -164 -147 -162
rect -153 -169 -147 -164
rect -153 -171 -150 -169
rect -148 -171 -147 -169
rect -153 -173 -147 -171
rect -153 -181 -149 -173
rect -137 -170 -99 -169
rect -137 -172 -103 -170
rect -101 -172 -99 -170
rect -137 -173 -99 -172
rect -153 -183 -152 -181
rect -150 -183 -149 -181
rect -104 -176 -99 -173
rect -129 -178 -114 -177
rect -129 -180 -125 -178
rect -123 -180 -118 -178
rect -116 -180 -114 -178
rect -129 -181 -114 -180
rect -104 -178 -96 -176
rect -104 -180 -99 -178
rect -97 -180 -96 -178
rect -173 -193 -165 -192
rect -254 -196 -252 -194
rect -250 -196 -249 -194
rect -254 -198 -249 -196
rect -191 -194 -165 -193
rect -191 -196 -174 -194
rect -172 -196 -168 -194
rect -166 -196 -165 -194
rect -191 -197 -165 -196
rect -153 -193 -149 -183
rect -120 -190 -116 -181
rect -104 -182 -96 -180
rect -73 -166 -68 -161
rect -73 -168 -72 -166
rect -70 -168 -68 -166
rect -73 -170 -68 -168
rect -153 -194 -131 -193
rect -153 -196 -150 -194
rect -148 -196 -131 -194
rect -153 -197 -131 -196
rect -72 -189 -68 -170
rect -72 -191 -71 -189
rect -69 -191 -68 -189
rect -72 -192 -68 -191
rect -73 -194 -68 -192
rect -73 -196 -72 -194
rect -70 -196 -68 -194
rect -73 -198 -68 -196
rect -258 -204 -64 -203
rect -284 -209 -64 -204
rect -285 -211 -64 -209
rect -285 -359 -279 -211
rect -49 -218 -42 -147
rect 137 -135 141 -103
rect 136 -137 141 -135
rect 136 -139 137 -137
rect 139 -139 141 -137
rect 136 -143 141 -139
rect 145 -107 151 -105
rect 225 -104 230 -102
rect 225 -106 226 -104
rect 228 -106 230 -104
rect 145 -109 148 -107
rect 150 -109 151 -107
rect 145 -114 151 -109
rect 145 -116 148 -114
rect 150 -116 151 -114
rect 145 -118 151 -116
rect 145 -138 149 -118
rect 161 -115 199 -114
rect 161 -117 187 -115
rect 189 -117 199 -115
rect 161 -118 199 -117
rect 194 -121 199 -118
rect 169 -123 184 -122
rect 169 -125 173 -123
rect 175 -125 180 -123
rect 182 -125 184 -123
rect 169 -126 184 -125
rect 194 -123 202 -121
rect 194 -125 199 -123
rect 201 -125 202 -123
rect 178 -132 182 -126
rect 194 -127 202 -125
rect 225 -111 230 -106
rect 225 -113 226 -111
rect 228 -113 230 -111
rect 225 -115 230 -113
rect 178 -134 179 -132
rect 181 -134 182 -132
rect 178 -135 182 -134
rect 145 -139 167 -138
rect 145 -141 148 -139
rect 150 -141 167 -139
rect 145 -142 167 -141
rect 226 -137 230 -115
rect 225 -139 230 -137
rect 225 -141 226 -139
rect 228 -141 230 -139
rect 225 -143 230 -141
rect 236 -102 249 -98
rect 325 -101 338 -98
rect 236 -104 241 -102
rect 236 -106 238 -104
rect 240 -106 241 -104
rect 325 -103 327 -101
rect 329 -102 338 -101
rect 365 -102 378 -98
rect 526 -102 539 -98
rect 566 -101 579 -98
rect 566 -102 575 -101
rect 236 -111 241 -106
rect 236 -113 238 -111
rect 240 -113 241 -111
rect 236 -115 241 -113
rect 236 -137 240 -115
rect 267 -115 305 -114
rect 267 -117 285 -115
rect 287 -117 305 -115
rect 267 -118 305 -117
rect 267 -121 272 -118
rect 264 -123 272 -121
rect 264 -125 265 -123
rect 267 -125 272 -123
rect 264 -127 272 -125
rect 282 -123 297 -122
rect 282 -125 284 -123
rect 286 -125 291 -123
rect 293 -125 297 -123
rect 282 -126 297 -125
rect 236 -139 241 -137
rect 284 -132 288 -126
rect 315 -107 321 -105
rect 315 -109 316 -107
rect 318 -109 321 -107
rect 315 -114 321 -109
rect 315 -116 316 -114
rect 318 -116 321 -114
rect 315 -118 321 -116
rect 284 -134 285 -132
rect 287 -134 288 -132
rect 284 -135 288 -134
rect 317 -138 321 -118
rect 236 -141 238 -139
rect 240 -141 241 -139
rect 236 -143 241 -141
rect 299 -139 321 -138
rect 299 -141 316 -139
rect 318 -141 321 -139
rect 299 -142 321 -141
rect 325 -107 329 -103
rect 365 -104 370 -102
rect 325 -109 326 -107
rect 328 -109 329 -107
rect 325 -135 329 -109
rect 349 -114 353 -105
rect 365 -106 367 -104
rect 369 -106 370 -104
rect 365 -111 370 -106
rect 365 -113 367 -111
rect 369 -113 370 -111
rect 340 -115 353 -114
rect 340 -117 341 -115
rect 343 -117 344 -115
rect 346 -117 353 -115
rect 340 -118 353 -117
rect 357 -114 361 -113
rect 357 -116 358 -114
rect 360 -116 361 -114
rect 357 -122 361 -116
rect 348 -123 361 -122
rect 348 -125 354 -123
rect 356 -125 361 -123
rect 348 -126 361 -125
rect 357 -127 361 -126
rect 365 -115 370 -113
rect 365 -123 369 -115
rect 365 -125 366 -123
rect 368 -125 369 -123
rect 396 -118 434 -114
rect 325 -137 330 -135
rect 325 -139 327 -137
rect 329 -139 330 -137
rect 325 -143 330 -139
rect 365 -137 369 -125
rect 396 -121 401 -118
rect 393 -123 401 -121
rect 393 -125 394 -123
rect 396 -125 398 -123
rect 400 -125 401 -123
rect 393 -127 401 -125
rect 411 -123 426 -122
rect 411 -125 413 -123
rect 415 -125 420 -123
rect 422 -125 426 -123
rect 411 -126 426 -125
rect 413 -128 414 -126
rect 416 -128 417 -126
rect 444 -107 450 -105
rect 444 -109 445 -107
rect 447 -109 450 -107
rect 444 -114 450 -109
rect 444 -116 445 -114
rect 447 -116 450 -114
rect 444 -118 450 -116
rect 365 -139 370 -137
rect 413 -135 417 -128
rect 446 -138 450 -118
rect 365 -141 367 -139
rect 369 -141 370 -139
rect 365 -143 370 -141
rect 428 -139 450 -138
rect 428 -141 445 -139
rect 447 -141 450 -139
rect 428 -142 450 -141
rect 454 -107 460 -105
rect 534 -104 539 -102
rect 534 -106 535 -104
rect 537 -106 539 -104
rect 454 -109 457 -107
rect 459 -109 460 -107
rect 454 -114 460 -109
rect 454 -116 457 -114
rect 459 -116 460 -114
rect 454 -118 460 -116
rect 454 -138 458 -118
rect 470 -118 508 -114
rect 503 -121 508 -118
rect 478 -123 493 -122
rect 478 -125 482 -123
rect 484 -125 489 -123
rect 491 -125 493 -123
rect 478 -126 493 -125
rect 503 -123 511 -121
rect 503 -125 505 -123
rect 507 -125 508 -123
rect 510 -125 511 -123
rect 487 -127 491 -126
rect 503 -127 511 -125
rect 487 -129 488 -127
rect 490 -129 491 -127
rect 487 -135 491 -129
rect 534 -111 539 -106
rect 534 -113 535 -111
rect 537 -113 539 -111
rect 534 -115 539 -113
rect 535 -123 539 -115
rect 535 -125 536 -123
rect 538 -125 539 -123
rect 454 -139 476 -138
rect 454 -141 457 -139
rect 459 -141 476 -139
rect 454 -142 476 -141
rect 535 -137 539 -125
rect 543 -114 547 -113
rect 543 -116 544 -114
rect 546 -116 547 -114
rect 543 -122 547 -116
rect 551 -114 555 -105
rect 577 -103 579 -101
rect 655 -102 668 -98
rect 747 -102 760 -98
rect 575 -105 579 -103
rect 551 -115 564 -114
rect 551 -117 558 -115
rect 560 -117 561 -115
rect 563 -117 564 -115
rect 551 -118 564 -117
rect 543 -123 556 -122
rect 543 -125 548 -123
rect 550 -125 556 -123
rect 543 -126 556 -125
rect 543 -127 547 -126
rect 575 -107 576 -105
rect 578 -107 579 -105
rect 534 -139 539 -137
rect 534 -141 535 -139
rect 537 -141 539 -139
rect 534 -143 539 -141
rect 575 -135 579 -107
rect 574 -137 579 -135
rect 574 -139 575 -137
rect 577 -139 579 -137
rect 574 -143 579 -139
rect 583 -107 589 -105
rect 663 -104 668 -102
rect 663 -106 664 -104
rect 666 -106 668 -104
rect 583 -109 586 -107
rect 588 -109 589 -107
rect 583 -114 589 -109
rect 583 -116 586 -114
rect 588 -116 589 -114
rect 583 -118 589 -116
rect 583 -138 587 -118
rect 599 -115 637 -114
rect 599 -117 623 -115
rect 625 -117 637 -115
rect 599 -118 637 -117
rect 632 -121 637 -118
rect 607 -123 622 -122
rect 607 -125 611 -123
rect 613 -125 618 -123
rect 620 -125 622 -123
rect 607 -126 622 -125
rect 632 -123 640 -121
rect 632 -125 637 -123
rect 639 -125 640 -123
rect 616 -132 620 -126
rect 632 -127 640 -125
rect 663 -111 668 -106
rect 663 -113 664 -111
rect 666 -113 668 -111
rect 663 -115 668 -113
rect 616 -134 617 -132
rect 619 -134 620 -132
rect 616 -135 620 -134
rect 583 -139 605 -138
rect 583 -141 586 -139
rect 588 -141 605 -139
rect 583 -142 605 -141
rect 664 -136 668 -115
rect 664 -137 665 -136
rect 663 -138 665 -137
rect 667 -138 668 -136
rect 663 -139 668 -138
rect 663 -141 664 -139
rect 666 -141 668 -139
rect 663 -143 668 -141
rect 675 -107 681 -105
rect 755 -104 760 -102
rect 755 -106 756 -104
rect 758 -106 760 -104
rect 675 -109 678 -107
rect 680 -109 681 -107
rect 675 -114 681 -109
rect 675 -116 678 -114
rect 680 -116 681 -114
rect 675 -118 681 -116
rect 675 -124 679 -118
rect 691 -115 729 -114
rect 691 -117 692 -115
rect 694 -117 729 -115
rect 691 -118 729 -117
rect 675 -126 676 -124
rect 678 -126 679 -124
rect 675 -138 679 -126
rect 724 -121 729 -118
rect 699 -123 713 -122
rect 699 -125 700 -123
rect 702 -125 703 -123
rect 705 -125 710 -123
rect 712 -125 713 -123
rect 699 -126 713 -125
rect 708 -127 713 -126
rect 724 -123 732 -121
rect 724 -125 729 -123
rect 731 -125 732 -123
rect 724 -127 732 -125
rect 708 -135 712 -127
rect 755 -111 760 -106
rect 755 -113 756 -111
rect 758 -113 760 -111
rect 755 -115 760 -113
rect 756 -123 760 -115
rect 756 -126 757 -123
rect 759 -126 760 -123
rect 675 -139 697 -138
rect 675 -141 678 -139
rect 680 -141 697 -139
rect 675 -142 697 -141
rect 756 -137 760 -126
rect 755 -139 760 -137
rect 755 -141 756 -139
rect 758 -141 760 -139
rect 755 -143 760 -141
rect 784 -148 790 31
rect 14 -149 794 -148
rect 14 -151 108 -149
rect 110 -151 136 -149
rect 138 -151 328 -149
rect 330 -151 356 -149
rect 358 -151 546 -149
rect 548 -151 574 -149
rect 576 -151 794 -149
rect 14 -156 794 -151
rect 636 -211 780 -208
rect 636 -213 638 -211
rect 640 -213 775 -211
rect 777 -213 780 -211
rect 636 -216 780 -213
rect -49 -223 569 -218
rect -49 -225 403 -223
rect 405 -225 417 -223
rect 419 -225 431 -223
rect 433 -225 446 -223
rect 448 -225 460 -223
rect 462 -225 474 -223
rect 476 -225 489 -223
rect 491 -225 503 -223
rect 505 -225 517 -223
rect 519 -225 532 -223
rect 534 -225 546 -223
rect 548 -225 560 -223
rect 562 -225 569 -223
rect -49 -226 569 -225
rect -49 -295 -42 -226
rect -256 -296 -42 -295
rect -256 -300 -43 -296
rect -256 -302 -249 -300
rect -247 -302 -235 -300
rect -233 -302 -221 -300
rect -219 -302 -206 -300
rect -204 -302 -192 -300
rect -190 -302 -178 -300
rect -176 -302 -163 -300
rect -161 -302 -149 -300
rect -147 -302 -135 -300
rect -133 -302 -120 -300
rect -118 -302 -106 -300
rect -104 -302 -92 -300
rect -90 -302 -43 -300
rect -256 -303 -43 -302
rect -252 -325 -248 -316
rect -252 -327 -250 -325
rect -252 -341 -248 -327
rect -237 -310 -224 -308
rect -237 -312 -233 -310
rect -231 -312 -224 -310
rect -237 -314 -224 -312
rect -237 -321 -231 -314
rect -209 -325 -205 -316
rect -209 -327 -207 -325
rect -252 -343 -251 -341
rect -249 -343 -248 -341
rect -252 -348 -248 -343
rect -252 -350 -250 -348
rect -248 -350 -240 -348
rect -252 -354 -240 -350
rect -220 -341 -216 -332
rect -229 -342 -216 -341
rect -229 -344 -224 -342
rect -222 -344 -216 -342
rect -229 -346 -216 -344
rect -209 -342 -205 -327
rect -194 -310 -186 -308
rect -194 -312 -190 -310
rect -188 -312 -186 -310
rect -194 -314 -186 -312
rect -194 -321 -188 -314
rect -166 -325 -162 -316
rect -166 -327 -164 -325
rect -209 -344 -208 -342
rect -206 -344 -205 -342
rect -209 -348 -205 -344
rect -209 -350 -207 -348
rect -205 -350 -197 -348
rect -209 -354 -197 -350
rect -177 -341 -173 -332
rect -186 -342 -173 -341
rect -186 -344 -181 -342
rect -179 -344 -173 -342
rect -186 -346 -173 -344
rect -166 -342 -162 -327
rect -151 -321 -145 -316
rect -123 -325 -119 -316
rect -123 -327 -121 -325
rect -166 -344 -165 -342
rect -163 -344 -162 -342
rect -166 -348 -162 -344
rect -166 -350 -164 -348
rect -162 -350 -154 -348
rect -166 -354 -154 -350
rect -134 -341 -130 -332
rect -143 -342 -130 -341
rect -143 -344 -138 -342
rect -136 -344 -130 -342
rect -143 -346 -130 -344
rect -123 -342 -119 -327
rect -108 -310 -95 -308
rect -108 -312 -104 -310
rect -102 -312 -95 -310
rect -108 -314 -95 -312
rect -108 -321 -102 -314
rect -123 -344 -122 -342
rect -120 -344 -119 -342
rect -123 -348 -119 -344
rect -123 -350 -121 -348
rect -119 -350 -111 -348
rect -123 -354 -111 -350
rect -91 -341 -87 -332
rect -100 -342 -87 -341
rect -100 -344 -95 -342
rect -93 -344 -87 -342
rect -100 -346 -87 -344
rect -285 -360 -83 -359
rect -285 -362 -249 -360
rect -247 -362 -239 -360
rect -237 -362 -206 -360
rect -204 -362 -196 -360
rect -194 -362 -163 -360
rect -161 -362 -153 -360
rect -151 -362 -120 -360
rect -118 -362 -110 -360
rect -108 -362 -83 -360
rect -285 -366 -83 -362
rect -285 -383 -279 -366
rect -256 -367 -83 -366
rect -68 -361 -63 -303
rect 367 -314 374 -226
rect 400 -248 404 -239
rect 400 -250 402 -248
rect 400 -264 404 -250
rect 415 -233 428 -231
rect 415 -235 419 -233
rect 421 -235 428 -233
rect 415 -237 428 -235
rect 415 -244 421 -237
rect 443 -248 447 -239
rect 443 -250 445 -248
rect 432 -257 436 -255
rect 432 -259 433 -257
rect 435 -259 436 -257
rect 400 -266 401 -264
rect 403 -266 404 -264
rect 400 -271 404 -266
rect 400 -273 402 -271
rect 404 -273 412 -271
rect 400 -277 412 -273
rect 432 -264 436 -259
rect 423 -265 436 -264
rect 423 -267 428 -265
rect 430 -267 436 -265
rect 423 -269 436 -267
rect 443 -265 447 -250
rect 458 -233 466 -231
rect 458 -235 462 -233
rect 464 -235 466 -233
rect 458 -237 466 -235
rect 458 -244 464 -237
rect 486 -248 490 -239
rect 486 -250 488 -248
rect 443 -267 444 -265
rect 446 -267 447 -265
rect 443 -271 447 -267
rect 443 -273 445 -271
rect 447 -273 455 -271
rect 443 -277 455 -273
rect 475 -264 479 -255
rect 466 -265 479 -264
rect 466 -267 471 -265
rect 473 -267 479 -265
rect 466 -269 479 -267
rect 486 -265 490 -250
rect 501 -244 507 -239
rect 529 -248 533 -239
rect 529 -250 531 -248
rect 486 -267 487 -265
rect 489 -267 490 -265
rect 486 -271 490 -267
rect 486 -273 488 -271
rect 490 -273 498 -271
rect 486 -277 498 -273
rect 518 -264 522 -255
rect 509 -265 522 -264
rect 509 -267 514 -265
rect 516 -267 522 -265
rect 509 -269 522 -267
rect 529 -271 533 -250
rect 544 -233 557 -231
rect 544 -235 548 -233
rect 550 -235 554 -233
rect 556 -235 557 -233
rect 544 -237 557 -235
rect 544 -244 550 -237
rect 529 -273 531 -271
rect 533 -273 541 -271
rect 529 -277 541 -273
rect 561 -264 565 -255
rect 552 -265 565 -264
rect 552 -267 557 -265
rect 559 -267 565 -265
rect 552 -269 565 -267
rect 396 -283 569 -282
rect 786 -283 794 -156
rect 396 -285 403 -283
rect 405 -285 413 -283
rect 415 -285 446 -283
rect 448 -285 456 -283
rect 458 -285 489 -283
rect 491 -285 499 -283
rect 501 -285 532 -283
rect 534 -285 542 -283
rect 544 -284 794 -283
rect 544 -285 793 -284
rect 396 -290 793 -285
rect 568 -291 793 -290
rect 590 -306 595 -303
rect 590 -308 591 -306
rect 593 -308 595 -306
rect 590 -309 595 -308
rect 367 -322 589 -314
rect 399 -332 412 -328
rect 572 -332 585 -328
rect 399 -334 404 -332
rect 399 -336 401 -334
rect 403 -336 404 -334
rect 399 -341 404 -336
rect 399 -343 401 -341
rect 403 -343 404 -341
rect 399 -345 404 -343
rect 399 -356 403 -345
rect 430 -345 468 -344
rect 430 -347 440 -345
rect 442 -347 468 -345
rect 430 -348 468 -347
rect 399 -358 400 -356
rect 402 -358 403 -356
rect -68 -362 18 -361
rect -286 -384 -279 -383
rect -68 -372 27 -362
rect -286 -456 -278 -384
rect -68 -391 -63 -372
rect -257 -399 -63 -391
rect -253 -409 -240 -405
rect -80 -409 -67 -405
rect -253 -411 -248 -409
rect -253 -413 -251 -411
rect -249 -413 -248 -411
rect -253 -418 -248 -413
rect -253 -420 -251 -418
rect -249 -420 -248 -418
rect -253 -422 -248 -420
rect -253 -432 -249 -422
rect -222 -422 -184 -421
rect -222 -424 -212 -422
rect -210 -424 -184 -422
rect -222 -425 -184 -424
rect -253 -434 -252 -432
rect -250 -434 -249 -432
rect -253 -444 -249 -434
rect -222 -428 -217 -425
rect -225 -430 -217 -428
rect -225 -432 -224 -430
rect -222 -432 -217 -430
rect -225 -434 -217 -432
rect -207 -430 -192 -429
rect -207 -432 -205 -430
rect -203 -432 -198 -430
rect -196 -432 -192 -430
rect -207 -433 -192 -432
rect -205 -434 -201 -433
rect -174 -414 -168 -412
rect -174 -416 -173 -414
rect -171 -416 -168 -414
rect -174 -421 -168 -416
rect -174 -423 -173 -421
rect -171 -423 -168 -421
rect -174 -425 -168 -423
rect -205 -436 -204 -434
rect -202 -436 -201 -434
rect -253 -446 -248 -444
rect -205 -442 -201 -436
rect -172 -443 -168 -425
rect -152 -414 -146 -412
rect -72 -411 -67 -409
rect -72 -413 -71 -411
rect -69 -413 -67 -411
rect -152 -416 -149 -414
rect -147 -416 -146 -414
rect -152 -421 -146 -416
rect -152 -423 -149 -421
rect -147 -423 -146 -421
rect -152 -425 -146 -423
rect -152 -433 -148 -425
rect -136 -422 -98 -421
rect -136 -424 -102 -422
rect -100 -424 -98 -422
rect -136 -425 -98 -424
rect -152 -435 -151 -433
rect -149 -435 -148 -433
rect -103 -428 -98 -425
rect -128 -430 -113 -429
rect -128 -432 -124 -430
rect -122 -432 -117 -430
rect -115 -432 -113 -430
rect -128 -433 -113 -432
rect -103 -430 -95 -428
rect -103 -432 -98 -430
rect -96 -432 -95 -430
rect -172 -445 -164 -443
rect -253 -448 -251 -446
rect -249 -448 -248 -446
rect -253 -450 -248 -448
rect -190 -446 -167 -445
rect -190 -448 -173 -446
rect -171 -447 -167 -446
rect -165 -447 -164 -445
rect -171 -448 -164 -447
rect -190 -449 -164 -448
rect -152 -445 -148 -435
rect -119 -442 -115 -433
rect -103 -434 -95 -432
rect -72 -418 -67 -413
rect -72 -420 -71 -418
rect -69 -420 -67 -418
rect -72 -422 -67 -420
rect -71 -433 -67 -422
rect -71 -435 -70 -433
rect -68 -435 -67 -433
rect -152 -446 -130 -445
rect -152 -448 -149 -446
rect -147 -448 -130 -446
rect -152 -449 -130 -448
rect -71 -444 -67 -435
rect -72 -446 -67 -444
rect -72 -448 -71 -446
rect -69 -448 -67 -446
rect -72 -450 -67 -448
rect -257 -456 -63 -455
rect -286 -463 -63 -456
rect 17 -459 27 -372
rect 399 -367 403 -358
rect 430 -351 435 -348
rect 427 -353 435 -351
rect 427 -355 428 -353
rect 430 -355 435 -353
rect 427 -357 435 -355
rect 445 -353 460 -352
rect 445 -355 447 -353
rect 449 -355 454 -353
rect 456 -355 460 -353
rect 445 -356 460 -355
rect 447 -357 451 -356
rect 478 -337 484 -335
rect 478 -339 479 -337
rect 481 -339 484 -337
rect 478 -344 484 -339
rect 478 -346 479 -344
rect 481 -346 484 -344
rect 478 -348 484 -346
rect 447 -359 448 -357
rect 450 -359 451 -357
rect 399 -369 404 -367
rect 447 -365 451 -359
rect 480 -367 484 -348
rect 500 -337 506 -335
rect 580 -334 585 -332
rect 580 -336 581 -334
rect 583 -336 585 -334
rect 500 -339 503 -337
rect 505 -339 506 -337
rect 500 -344 506 -339
rect 500 -346 503 -344
rect 505 -346 506 -344
rect 500 -348 506 -346
rect 500 -356 504 -348
rect 516 -345 554 -344
rect 516 -347 550 -345
rect 552 -347 554 -345
rect 516 -348 554 -347
rect 500 -358 501 -356
rect 503 -358 504 -356
rect 549 -351 554 -348
rect 524 -353 539 -352
rect 524 -355 528 -353
rect 530 -355 535 -353
rect 537 -355 539 -353
rect 524 -356 539 -355
rect 549 -353 557 -351
rect 549 -355 554 -353
rect 556 -355 557 -353
rect 480 -368 487 -367
rect 399 -371 401 -369
rect 403 -371 404 -369
rect 399 -373 404 -371
rect 462 -369 487 -368
rect 462 -371 479 -369
rect 481 -371 484 -369
rect 486 -371 487 -369
rect 462 -372 487 -371
rect 500 -368 504 -358
rect 533 -365 537 -356
rect 549 -357 557 -355
rect 580 -341 585 -336
rect 580 -343 581 -341
rect 583 -343 585 -341
rect 580 -345 585 -343
rect 500 -369 522 -368
rect 500 -371 503 -369
rect 505 -371 522 -369
rect 500 -372 522 -371
rect 581 -367 585 -345
rect 580 -369 585 -367
rect 580 -371 581 -369
rect 583 -371 585 -369
rect 580 -373 585 -371
rect 624 -378 629 -291
rect 395 -382 629 -378
rect 395 -384 411 -382
rect 413 -384 629 -382
rect 395 -385 629 -384
rect 395 -386 589 -385
rect -286 -668 -278 -463
rect -15 -468 27 -459
rect -16 -469 27 -468
rect -16 -470 767 -469
rect -16 -603 -5 -470
rect 16 -474 767 -470
rect 16 -476 138 -474
rect 140 -476 330 -474
rect 332 -476 576 -474
rect 578 -476 767 -474
rect 16 -477 767 -476
rect 90 -487 103 -483
rect 130 -486 143 -483
rect 130 -487 139 -486
rect 18 -492 24 -490
rect 98 -489 103 -487
rect 98 -491 99 -489
rect 101 -491 103 -489
rect 18 -494 21 -492
rect 23 -494 24 -492
rect 18 -499 24 -494
rect 18 -501 21 -499
rect 23 -501 24 -499
rect 18 -503 24 -501
rect 18 -523 22 -503
rect 34 -503 72 -499
rect 67 -506 72 -503
rect 42 -508 57 -507
rect 42 -510 46 -508
rect 48 -510 53 -508
rect 55 -510 57 -508
rect 42 -511 57 -510
rect 67 -508 75 -506
rect 67 -510 68 -508
rect 70 -510 72 -508
rect 74 -510 75 -508
rect 18 -524 40 -523
rect 18 -526 21 -524
rect 23 -526 40 -524
rect 18 -527 40 -526
rect 51 -533 55 -511
rect 67 -512 75 -510
rect 98 -496 103 -491
rect 98 -498 99 -496
rect 101 -498 103 -496
rect 98 -500 103 -498
rect 99 -508 103 -500
rect 99 -510 100 -508
rect 102 -510 103 -508
rect 99 -522 103 -510
rect 107 -499 111 -498
rect 107 -501 108 -499
rect 110 -501 111 -499
rect 107 -507 111 -501
rect 115 -499 119 -490
rect 141 -488 143 -486
rect 219 -487 232 -483
rect 115 -500 128 -499
rect 115 -502 122 -500
rect 124 -502 125 -500
rect 127 -502 128 -500
rect 115 -503 128 -502
rect 107 -508 120 -507
rect 107 -510 112 -508
rect 114 -510 120 -508
rect 107 -511 120 -510
rect 107 -512 111 -511
rect 98 -524 103 -522
rect 98 -526 99 -524
rect 101 -526 103 -524
rect 98 -528 103 -526
rect 139 -520 143 -488
rect 138 -522 143 -520
rect 138 -524 139 -522
rect 141 -524 143 -522
rect 138 -528 143 -524
rect 147 -492 153 -490
rect 227 -489 232 -487
rect 227 -491 228 -489
rect 230 -491 232 -489
rect 147 -494 150 -492
rect 152 -494 153 -492
rect 147 -499 153 -494
rect 147 -501 150 -499
rect 152 -501 153 -499
rect 147 -503 153 -501
rect 147 -523 151 -503
rect 163 -500 201 -499
rect 163 -502 189 -500
rect 191 -502 201 -500
rect 163 -503 201 -502
rect 196 -506 201 -503
rect 171 -508 186 -507
rect 171 -510 175 -508
rect 177 -510 182 -508
rect 184 -510 186 -508
rect 171 -511 186 -510
rect 196 -508 204 -506
rect 196 -510 201 -508
rect 203 -510 204 -508
rect 180 -517 184 -511
rect 196 -512 204 -510
rect 227 -496 232 -491
rect 227 -498 228 -496
rect 230 -498 232 -496
rect 227 -500 232 -498
rect 180 -519 181 -517
rect 183 -519 184 -517
rect 180 -520 184 -519
rect 147 -524 169 -523
rect 147 -526 150 -524
rect 152 -526 169 -524
rect 147 -527 169 -526
rect 228 -522 232 -500
rect 227 -524 232 -522
rect 227 -526 228 -524
rect 230 -526 232 -524
rect 227 -528 232 -526
rect 238 -487 251 -483
rect 327 -486 340 -483
rect 238 -489 243 -487
rect 238 -491 240 -489
rect 242 -491 243 -489
rect 327 -488 329 -486
rect 331 -487 340 -486
rect 367 -487 380 -483
rect 528 -487 541 -483
rect 568 -486 581 -483
rect 568 -487 577 -486
rect 238 -496 243 -491
rect 238 -498 240 -496
rect 242 -498 243 -496
rect 238 -500 243 -498
rect 238 -522 242 -500
rect 269 -500 307 -499
rect 269 -502 287 -500
rect 289 -502 307 -500
rect 269 -503 307 -502
rect 269 -506 274 -503
rect 266 -508 274 -506
rect 266 -510 267 -508
rect 269 -510 274 -508
rect 266 -512 274 -510
rect 284 -508 299 -507
rect 284 -510 286 -508
rect 288 -510 293 -508
rect 295 -510 299 -508
rect 284 -511 299 -510
rect 238 -524 243 -522
rect 286 -517 290 -511
rect 317 -492 323 -490
rect 317 -494 318 -492
rect 320 -494 323 -492
rect 317 -499 323 -494
rect 317 -501 318 -499
rect 320 -501 323 -499
rect 317 -503 323 -501
rect 286 -519 287 -517
rect 289 -519 290 -517
rect 286 -520 290 -519
rect 319 -523 323 -503
rect 238 -526 240 -524
rect 242 -526 243 -524
rect 238 -528 243 -526
rect 301 -524 323 -523
rect 301 -526 318 -524
rect 320 -526 323 -524
rect 301 -527 323 -526
rect 327 -492 331 -488
rect 367 -489 372 -487
rect 327 -494 328 -492
rect 330 -494 331 -492
rect 327 -520 331 -494
rect 351 -499 355 -490
rect 367 -491 369 -489
rect 371 -491 372 -489
rect 367 -496 372 -491
rect 367 -498 369 -496
rect 371 -498 372 -496
rect 342 -500 355 -499
rect 342 -502 343 -500
rect 345 -502 346 -500
rect 348 -502 355 -500
rect 342 -503 355 -502
rect 359 -499 363 -498
rect 359 -501 360 -499
rect 362 -501 363 -499
rect 359 -507 363 -501
rect 350 -508 363 -507
rect 350 -510 356 -508
rect 358 -510 363 -508
rect 350 -511 363 -510
rect 359 -512 363 -511
rect 367 -500 372 -498
rect 367 -508 371 -500
rect 367 -510 368 -508
rect 370 -510 371 -508
rect 398 -503 436 -499
rect 327 -522 332 -520
rect 327 -524 329 -522
rect 331 -524 332 -522
rect 327 -528 332 -524
rect 367 -522 371 -510
rect 398 -506 403 -503
rect 395 -508 403 -506
rect 395 -510 396 -508
rect 398 -510 400 -508
rect 402 -510 403 -508
rect 395 -512 403 -510
rect 413 -508 428 -507
rect 413 -510 415 -508
rect 417 -510 422 -508
rect 424 -510 428 -508
rect 413 -511 428 -510
rect 367 -524 372 -522
rect 415 -516 419 -511
rect 446 -492 452 -490
rect 446 -494 447 -492
rect 449 -494 452 -492
rect 446 -499 452 -494
rect 446 -501 447 -499
rect 449 -501 452 -499
rect 446 -503 452 -501
rect 415 -518 416 -516
rect 418 -518 419 -516
rect 415 -520 419 -518
rect 448 -523 452 -503
rect 367 -526 369 -524
rect 371 -526 372 -524
rect 367 -528 372 -526
rect 430 -524 452 -523
rect 430 -526 447 -524
rect 449 -526 452 -524
rect 430 -527 452 -526
rect 456 -492 462 -490
rect 536 -489 541 -487
rect 536 -491 537 -489
rect 539 -491 541 -489
rect 456 -494 459 -492
rect 461 -494 462 -492
rect 456 -499 462 -494
rect 456 -501 459 -499
rect 461 -501 462 -499
rect 456 -503 462 -501
rect 456 -523 460 -503
rect 472 -503 510 -499
rect 505 -506 510 -503
rect 480 -508 495 -507
rect 480 -510 484 -508
rect 486 -510 491 -508
rect 493 -510 495 -508
rect 480 -511 495 -510
rect 505 -508 513 -506
rect 505 -510 506 -508
rect 508 -510 510 -508
rect 512 -510 513 -508
rect 489 -517 493 -511
rect 505 -512 513 -510
rect 536 -496 541 -491
rect 536 -498 537 -496
rect 539 -498 541 -496
rect 536 -500 541 -498
rect 537 -508 541 -500
rect 537 -510 538 -508
rect 540 -510 541 -508
rect 489 -519 490 -517
rect 492 -519 493 -517
rect 489 -520 493 -519
rect 456 -524 478 -523
rect 456 -526 459 -524
rect 461 -526 478 -524
rect 456 -527 478 -526
rect 537 -522 541 -510
rect 545 -499 549 -498
rect 545 -501 546 -499
rect 548 -501 549 -499
rect 545 -507 549 -501
rect 553 -499 557 -490
rect 579 -488 581 -486
rect 657 -487 670 -483
rect 749 -487 762 -483
rect 577 -490 581 -488
rect 553 -500 566 -499
rect 553 -502 560 -500
rect 562 -502 563 -500
rect 565 -502 566 -500
rect 553 -503 566 -502
rect 545 -508 558 -507
rect 545 -510 550 -508
rect 552 -510 558 -508
rect 545 -511 558 -510
rect 545 -512 549 -511
rect 577 -492 578 -490
rect 580 -492 581 -490
rect 536 -524 541 -522
rect 536 -526 537 -524
rect 539 -526 541 -524
rect 536 -528 541 -526
rect 577 -520 581 -492
rect 576 -522 581 -520
rect 576 -524 577 -522
rect 579 -524 581 -522
rect 576 -528 581 -524
rect 585 -492 591 -490
rect 665 -489 670 -487
rect 665 -491 666 -489
rect 668 -491 670 -489
rect 585 -494 588 -492
rect 590 -494 591 -492
rect 585 -499 591 -494
rect 585 -501 588 -499
rect 590 -501 591 -499
rect 585 -503 591 -501
rect 585 -523 589 -503
rect 601 -500 639 -499
rect 601 -502 625 -500
rect 627 -502 639 -500
rect 601 -503 639 -502
rect 634 -506 639 -503
rect 609 -508 624 -507
rect 609 -510 613 -508
rect 615 -510 620 -508
rect 622 -510 624 -508
rect 609 -511 624 -510
rect 634 -508 642 -506
rect 634 -510 639 -508
rect 641 -510 642 -508
rect 618 -517 622 -511
rect 634 -512 642 -510
rect 665 -496 670 -491
rect 665 -498 666 -496
rect 668 -498 670 -496
rect 665 -500 670 -498
rect 618 -519 619 -517
rect 621 -519 622 -517
rect 618 -520 622 -519
rect 585 -524 607 -523
rect 585 -526 588 -524
rect 590 -526 607 -524
rect 585 -527 607 -526
rect 666 -522 670 -500
rect 665 -524 670 -522
rect 665 -526 666 -524
rect 668 -526 670 -524
rect 665 -528 670 -526
rect 677 -492 683 -490
rect 757 -489 762 -487
rect 757 -491 758 -489
rect 760 -491 762 -489
rect 677 -494 680 -492
rect 682 -494 683 -492
rect 677 -499 683 -494
rect 677 -501 680 -499
rect 682 -501 683 -499
rect 677 -503 683 -501
rect 677 -509 681 -503
rect 693 -500 731 -499
rect 693 -502 718 -500
rect 720 -502 731 -500
rect 693 -503 731 -502
rect 677 -511 678 -509
rect 680 -511 681 -509
rect 677 -523 681 -511
rect 726 -506 731 -503
rect 701 -508 716 -507
rect 701 -510 702 -508
rect 704 -510 705 -508
rect 707 -510 712 -508
rect 714 -510 716 -508
rect 701 -511 716 -510
rect 726 -508 734 -506
rect 726 -510 731 -508
rect 733 -510 734 -508
rect 710 -520 714 -511
rect 726 -512 734 -510
rect 757 -496 762 -491
rect 757 -498 758 -496
rect 760 -498 762 -496
rect 757 -500 762 -498
rect 677 -524 699 -523
rect 677 -526 680 -524
rect 682 -526 699 -524
rect 677 -527 699 -526
rect 758 -522 762 -500
rect 757 -524 762 -522
rect 757 -526 758 -524
rect 760 -526 762 -524
rect 757 -528 762 -526
rect 786 -533 793 -291
rect 16 -534 794 -533
rect 16 -536 110 -534
rect 112 -536 138 -534
rect 140 -536 330 -534
rect 332 -536 358 -534
rect 360 -536 548 -534
rect 550 -536 576 -534
rect 578 -536 794 -534
rect 16 -541 794 -536
rect -251 -608 500 -603
rect -251 -610 -129 -608
rect -127 -610 63 -608
rect 65 -610 309 -608
rect 311 -610 500 -608
rect -251 -611 500 -610
rect -177 -621 -164 -617
rect -137 -620 -124 -617
rect -137 -621 -128 -620
rect -249 -626 -243 -624
rect -169 -623 -164 -621
rect -169 -625 -168 -623
rect -166 -625 -164 -623
rect -249 -628 -246 -626
rect -244 -628 -243 -626
rect -249 -633 -243 -628
rect -249 -635 -246 -633
rect -244 -635 -243 -633
rect -249 -637 -243 -635
rect -249 -657 -245 -637
rect -233 -637 -195 -633
rect -200 -640 -195 -637
rect -225 -642 -210 -641
rect -225 -644 -221 -642
rect -219 -644 -214 -642
rect -212 -644 -210 -642
rect -225 -645 -210 -644
rect -200 -642 -192 -640
rect -200 -644 -199 -642
rect -197 -644 -195 -642
rect -193 -644 -192 -642
rect -216 -651 -212 -645
rect -200 -646 -192 -644
rect -169 -630 -164 -625
rect -169 -632 -168 -630
rect -166 -632 -164 -630
rect -169 -634 -164 -632
rect -168 -642 -164 -634
rect -168 -644 -167 -642
rect -165 -644 -164 -642
rect -216 -653 -215 -651
rect -213 -653 -212 -651
rect -216 -654 -212 -653
rect -249 -658 -227 -657
rect -249 -660 -246 -658
rect -244 -660 -227 -658
rect -249 -661 -227 -660
rect -168 -656 -164 -644
rect -160 -633 -156 -632
rect -160 -635 -159 -633
rect -157 -635 -156 -633
rect -160 -641 -156 -635
rect -152 -633 -148 -624
rect -126 -622 -124 -620
rect -48 -621 -35 -617
rect -152 -634 -139 -633
rect -152 -636 -145 -634
rect -143 -636 -142 -634
rect -140 -636 -139 -634
rect -152 -637 -139 -636
rect -160 -642 -147 -641
rect -160 -644 -155 -642
rect -153 -644 -147 -642
rect -160 -645 -147 -644
rect -160 -646 -156 -645
rect -169 -658 -164 -656
rect -169 -660 -168 -658
rect -166 -660 -164 -658
rect -169 -662 -164 -660
rect -128 -654 -124 -622
rect -129 -656 -124 -654
rect -129 -658 -128 -656
rect -126 -658 -124 -656
rect -129 -662 -124 -658
rect -120 -626 -114 -624
rect -40 -623 -35 -621
rect -40 -625 -39 -623
rect -37 -625 -35 -623
rect -120 -628 -117 -626
rect -115 -628 -114 -626
rect -120 -633 -114 -628
rect -120 -635 -117 -633
rect -115 -635 -114 -633
rect -120 -637 -114 -635
rect -120 -657 -116 -637
rect -104 -634 -66 -633
rect -104 -636 -78 -634
rect -76 -636 -66 -634
rect -104 -637 -66 -636
rect -71 -640 -66 -637
rect -96 -642 -81 -641
rect -96 -644 -92 -642
rect -90 -644 -85 -642
rect -83 -644 -81 -642
rect -96 -645 -81 -644
rect -71 -642 -63 -640
rect -71 -644 -66 -642
rect -64 -644 -63 -642
rect -87 -651 -83 -645
rect -71 -646 -63 -644
rect -40 -630 -35 -625
rect -40 -632 -39 -630
rect -37 -632 -35 -630
rect -40 -634 -35 -632
rect -87 -653 -86 -651
rect -84 -653 -83 -651
rect -87 -654 -83 -653
rect -120 -658 -98 -657
rect -120 -660 -117 -658
rect -115 -660 -98 -658
rect -120 -661 -98 -660
rect -39 -656 -35 -634
rect -40 -658 -35 -656
rect -40 -660 -39 -658
rect -37 -660 -35 -658
rect -40 -662 -35 -660
rect -29 -621 -16 -617
rect 60 -620 73 -617
rect -29 -623 -24 -621
rect -29 -625 -27 -623
rect -25 -625 -24 -623
rect 60 -622 62 -620
rect 64 -621 73 -620
rect 100 -621 113 -617
rect 261 -621 274 -617
rect 301 -620 314 -617
rect 301 -621 310 -620
rect -29 -630 -24 -625
rect -29 -632 -27 -630
rect -25 -632 -24 -630
rect -29 -634 -24 -632
rect -29 -656 -25 -634
rect 2 -634 40 -633
rect 2 -636 20 -634
rect 22 -636 40 -634
rect 2 -637 40 -636
rect 2 -640 7 -637
rect -1 -642 7 -640
rect -1 -644 0 -642
rect 2 -644 7 -642
rect -1 -646 7 -644
rect 17 -642 32 -641
rect 17 -644 19 -642
rect 21 -644 26 -642
rect 28 -644 32 -642
rect 17 -645 32 -644
rect -29 -658 -24 -656
rect 19 -651 23 -645
rect 50 -626 56 -624
rect 50 -628 51 -626
rect 53 -628 56 -626
rect 50 -633 56 -628
rect 50 -635 51 -633
rect 53 -635 56 -633
rect 50 -637 56 -635
rect 19 -653 20 -651
rect 22 -653 23 -651
rect 19 -654 23 -653
rect 52 -657 56 -637
rect -29 -660 -27 -658
rect -25 -660 -24 -658
rect -29 -662 -24 -660
rect 34 -658 56 -657
rect 34 -660 51 -658
rect 53 -660 56 -658
rect 34 -661 56 -660
rect 60 -626 64 -622
rect 100 -623 105 -621
rect 60 -628 61 -626
rect 63 -628 64 -626
rect 60 -654 64 -628
rect 84 -633 88 -624
rect 100 -625 102 -623
rect 104 -625 105 -623
rect 100 -630 105 -625
rect 100 -632 102 -630
rect 104 -632 105 -630
rect 75 -634 88 -633
rect 75 -636 76 -634
rect 78 -636 79 -634
rect 81 -636 88 -634
rect 75 -637 88 -636
rect 92 -633 96 -632
rect 92 -635 93 -633
rect 95 -635 96 -633
rect 92 -641 96 -635
rect 83 -642 96 -641
rect 83 -644 89 -642
rect 91 -644 96 -642
rect 83 -645 96 -644
rect 92 -646 96 -645
rect 100 -634 105 -632
rect 100 -642 104 -634
rect 100 -644 101 -642
rect 103 -644 104 -642
rect 131 -637 169 -633
rect 60 -656 65 -654
rect 60 -658 62 -656
rect 64 -658 65 -656
rect 60 -662 65 -658
rect 100 -656 104 -644
rect 131 -640 136 -637
rect 128 -642 136 -640
rect 128 -644 129 -642
rect 131 -644 136 -642
rect 128 -646 136 -644
rect 146 -642 161 -641
rect 146 -644 148 -642
rect 150 -644 155 -642
rect 157 -644 161 -642
rect 146 -645 161 -644
rect 100 -658 105 -656
rect 148 -651 152 -645
rect 179 -626 185 -624
rect 179 -628 180 -626
rect 182 -628 185 -626
rect 179 -633 185 -628
rect 179 -635 180 -633
rect 182 -635 185 -633
rect 179 -637 185 -635
rect 148 -653 149 -651
rect 151 -653 152 -651
rect 148 -654 152 -653
rect 181 -657 185 -637
rect 100 -660 102 -658
rect 104 -660 105 -658
rect 100 -662 105 -660
rect 163 -658 185 -657
rect 163 -660 180 -658
rect 182 -660 185 -658
rect 163 -661 185 -660
rect 189 -626 195 -624
rect 269 -623 274 -621
rect 269 -625 270 -623
rect 272 -625 274 -623
rect 189 -628 192 -626
rect 194 -628 195 -626
rect 189 -633 195 -628
rect 189 -635 192 -633
rect 194 -635 195 -633
rect 189 -637 195 -635
rect 189 -657 193 -637
rect 205 -637 243 -633
rect 238 -640 243 -637
rect 213 -642 228 -641
rect 213 -644 217 -642
rect 219 -644 224 -642
rect 226 -644 228 -642
rect 213 -645 228 -644
rect 238 -642 246 -640
rect 238 -644 240 -642
rect 242 -644 243 -642
rect 245 -644 246 -642
rect 222 -651 226 -645
rect 238 -646 246 -644
rect 269 -630 274 -625
rect 269 -632 270 -630
rect 272 -632 274 -630
rect 269 -634 274 -632
rect 270 -642 274 -634
rect 270 -644 271 -642
rect 273 -644 274 -642
rect 222 -653 223 -651
rect 225 -653 226 -651
rect 222 -654 226 -653
rect 189 -658 211 -657
rect 189 -660 192 -658
rect 194 -660 211 -658
rect 189 -661 211 -660
rect 270 -656 274 -644
rect 278 -633 282 -632
rect 278 -635 279 -633
rect 281 -635 282 -633
rect 278 -641 282 -635
rect 286 -633 290 -624
rect 312 -622 314 -620
rect 390 -621 403 -617
rect 482 -621 495 -617
rect 310 -624 314 -622
rect 286 -634 299 -633
rect 286 -636 293 -634
rect 295 -636 296 -634
rect 298 -636 299 -634
rect 286 -637 299 -636
rect 278 -642 291 -641
rect 278 -644 283 -642
rect 285 -644 291 -642
rect 278 -645 291 -644
rect 278 -646 282 -645
rect 310 -626 311 -624
rect 313 -626 314 -624
rect 269 -658 274 -656
rect 269 -660 270 -658
rect 272 -660 274 -658
rect 269 -662 274 -660
rect 310 -654 314 -626
rect 309 -656 314 -654
rect 309 -658 310 -656
rect 312 -658 314 -656
rect 309 -662 314 -658
rect 318 -626 324 -624
rect 398 -623 403 -621
rect 398 -625 399 -623
rect 401 -625 403 -623
rect 318 -628 321 -626
rect 323 -628 324 -626
rect 318 -633 324 -628
rect 318 -635 321 -633
rect 323 -635 324 -633
rect 318 -637 324 -635
rect 318 -657 322 -637
rect 334 -634 372 -633
rect 334 -636 358 -634
rect 360 -636 372 -634
rect 334 -637 372 -636
rect 367 -640 372 -637
rect 342 -642 357 -641
rect 342 -644 346 -642
rect 348 -644 353 -642
rect 355 -644 357 -642
rect 342 -645 357 -644
rect 367 -642 375 -640
rect 367 -644 372 -642
rect 374 -644 375 -642
rect 351 -651 355 -645
rect 367 -646 375 -644
rect 398 -630 403 -625
rect 398 -632 399 -630
rect 401 -632 403 -630
rect 398 -634 403 -632
rect 351 -653 352 -651
rect 354 -653 355 -651
rect 351 -654 355 -653
rect 318 -658 340 -657
rect 318 -660 321 -658
rect 323 -660 340 -658
rect 318 -661 340 -660
rect 399 -656 403 -634
rect 398 -658 403 -656
rect 398 -660 399 -658
rect 401 -660 403 -658
rect 398 -662 403 -660
rect 410 -626 416 -624
rect 490 -623 495 -621
rect 490 -625 491 -623
rect 493 -625 495 -623
rect 410 -628 413 -626
rect 415 -628 416 -626
rect 410 -633 416 -628
rect 410 -635 413 -633
rect 415 -635 416 -633
rect 410 -637 416 -635
rect 410 -643 414 -637
rect 426 -634 464 -633
rect 426 -636 453 -634
rect 455 -636 464 -634
rect 426 -637 464 -636
rect 410 -645 411 -643
rect 413 -645 414 -643
rect 410 -657 414 -645
rect 459 -640 464 -637
rect 434 -642 449 -641
rect 434 -644 438 -642
rect 440 -644 445 -642
rect 447 -644 449 -642
rect 434 -645 449 -644
rect 459 -642 467 -640
rect 459 -644 464 -642
rect 466 -644 467 -642
rect 443 -654 447 -645
rect 459 -646 467 -644
rect 490 -630 495 -625
rect 490 -632 491 -630
rect 493 -632 495 -630
rect 490 -634 495 -632
rect 410 -658 432 -657
rect 410 -660 413 -658
rect 415 -660 432 -658
rect 410 -661 432 -660
rect 491 -656 495 -634
rect 490 -658 495 -656
rect 490 -660 491 -658
rect 493 -660 495 -658
rect 490 -662 495 -660
rect -251 -668 500 -667
rect -286 -670 -157 -668
rect -155 -670 -129 -668
rect -127 -670 63 -668
rect 65 -670 91 -668
rect 93 -669 281 -668
rect 93 -670 149 -669
rect -286 -671 149 -670
rect 151 -670 281 -669
rect 283 -670 309 -668
rect 311 -670 500 -668
rect 151 -671 500 -670
rect -286 -675 500 -671
rect 308 -680 324 -675
rect 308 -738 325 -680
rect 680 -738 697 -541
rect 767 -542 794 -541
rect -58 -739 800 -738
rect -336 -781 874 -739
<< alu2 >>
rect 100 210 419 214
rect 100 201 104 210
rect -33 199 104 201
rect -33 197 -31 199
rect -29 197 104 199
rect -33 196 104 197
rect 413 184 419 210
rect 413 182 415 184
rect 417 182 419 184
rect 413 180 419 182
rect 258 153 271 154
rect 258 151 268 153
rect 270 151 271 153
rect 258 150 271 151
rect 304 152 314 153
rect 304 150 311 152
rect 313 150 314 152
rect 258 114 263 150
rect 304 149 314 150
rect 347 152 357 153
rect 347 150 354 152
rect 356 150 357 152
rect 347 149 357 150
rect 304 123 309 149
rect 304 118 340 123
rect 258 109 311 114
rect 306 72 311 109
rect 333 111 340 118
rect 347 121 352 149
rect 396 143 703 146
rect 396 141 398 143
rect 400 141 703 143
rect 396 140 703 141
rect 347 117 421 121
rect 333 105 401 111
rect 306 70 307 72
rect 309 70 311 72
rect 306 69 311 70
rect 393 64 399 105
rect 415 72 421 117
rect 415 70 417 72
rect 419 70 421 72
rect 415 69 421 70
rect 393 62 395 64
rect 397 62 399 64
rect 314 61 371 62
rect 314 60 368 61
rect 314 58 315 60
rect 317 59 368 60
rect 370 59 371 61
rect 393 60 399 62
rect 317 58 371 59
rect 314 57 371 58
rect 251 54 270 56
rect 251 52 267 54
rect 269 52 270 54
rect 448 55 500 57
rect 448 53 449 55
rect 451 53 495 55
rect 497 53 500 55
rect 251 51 270 52
rect 351 52 355 53
rect 448 52 500 53
rect 251 7 257 51
rect 251 5 253 7
rect 255 5 257 7
rect 251 3 257 5
rect 351 50 352 52
rect 354 50 355 52
rect -96 -13 344 -8
rect 351 -9 355 50
rect 351 -11 352 -9
rect 354 -11 355 -9
rect 351 -13 355 -11
rect 687 -10 691 -9
rect 687 -12 688 -10
rect 690 -12 691 -10
rect -96 -30 -92 -13
rect 340 -17 344 -13
rect 687 -17 691 -12
rect 340 -21 691 -17
rect -79 -25 -74 -22
rect -229 -36 -92 -30
rect -80 -27 659 -25
rect -80 -29 654 -27
rect 656 -29 659 -27
rect -80 -32 659 -29
rect -229 -58 -225 -36
rect -79 -56 -74 -32
rect -229 -60 -228 -58
rect -226 -60 -225 -58
rect -100 -57 -74 -56
rect -100 -59 -99 -57
rect -97 -59 -74 -57
rect -100 -60 -74 -59
rect -229 -62 -225 -60
rect -124 -66 695 -64
rect -124 -68 -123 -66
rect -121 -68 695 -66
rect -124 -70 695 -68
rect -262 -89 -249 -88
rect -262 -91 -252 -89
rect -250 -91 -249 -89
rect -262 -92 -249 -91
rect -216 -90 -206 -89
rect -216 -92 -209 -90
rect -207 -92 -206 -90
rect -262 -128 -257 -92
rect -216 -93 -206 -92
rect -173 -90 -163 -89
rect -173 -92 -166 -90
rect -164 -92 -163 -90
rect -173 -93 -163 -92
rect -216 -119 -211 -93
rect -216 -124 -180 -119
rect -262 -133 -209 -128
rect -214 -170 -209 -133
rect -187 -131 -180 -124
rect -173 -121 -168 -93
rect 128 -99 144 -98
rect 128 -101 129 -99
rect 131 -101 141 -99
rect 143 -101 144 -99
rect 128 -102 144 -101
rect 186 -102 329 -97
rect 18 -114 109 -113
rect 145 -114 151 -113
rect 18 -116 19 -114
rect 21 -116 106 -114
rect 108 -116 109 -114
rect 18 -117 109 -116
rect 122 -115 148 -114
rect 122 -117 123 -115
rect 125 -116 148 -115
rect 150 -116 151 -114
rect 125 -117 151 -116
rect 122 -118 151 -117
rect 186 -115 190 -102
rect 186 -117 187 -115
rect 189 -117 190 -115
rect 186 -118 190 -117
rect 284 -107 288 -106
rect 284 -109 285 -107
rect 287 -109 288 -107
rect 284 -115 288 -109
rect 325 -107 329 -102
rect 563 -102 579 -100
rect 563 -104 564 -102
rect 566 -104 579 -102
rect 563 -105 579 -104
rect 325 -109 326 -107
rect 328 -109 329 -107
rect 575 -107 576 -105
rect 578 -107 579 -105
rect 575 -109 579 -107
rect 622 -101 680 -95
rect 325 -110 329 -109
rect 284 -117 285 -115
rect 287 -117 288 -115
rect 284 -118 288 -117
rect 315 -114 321 -113
rect 357 -114 448 -113
rect 315 -116 316 -114
rect 318 -115 344 -114
rect 318 -116 341 -115
rect 315 -117 341 -116
rect 343 -117 344 -115
rect 357 -116 358 -114
rect 360 -116 445 -114
rect 447 -116 448 -114
rect 357 -117 448 -116
rect 456 -114 547 -113
rect 583 -114 589 -113
rect 456 -116 457 -114
rect 459 -116 544 -114
rect 546 -116 547 -114
rect 456 -117 547 -116
rect 560 -115 586 -114
rect 560 -117 561 -115
rect 563 -116 586 -115
rect 588 -116 589 -114
rect 563 -117 589 -116
rect 315 -118 344 -117
rect 560 -118 589 -117
rect 622 -115 627 -101
rect 622 -117 623 -115
rect 625 -117 627 -115
rect 622 -118 627 -117
rect -173 -125 -99 -121
rect -187 -137 -119 -131
rect -214 -172 -213 -170
rect -211 -172 -209 -170
rect -214 -173 -209 -172
rect -127 -178 -121 -137
rect -105 -170 -99 -125
rect 65 -123 70 -121
rect 65 -125 66 -123
rect 68 -125 70 -123
rect 49 -132 59 -131
rect 49 -134 50 -132
rect 52 -134 56 -132
rect 58 -134 59 -132
rect 49 -135 59 -134
rect -105 -172 -103 -170
rect -101 -172 -99 -170
rect -105 -173 -99 -172
rect -265 -180 -250 -178
rect -127 -180 -125 -178
rect -123 -180 -121 -178
rect -265 -182 -253 -180
rect -251 -182 -250 -180
rect -265 -183 -250 -182
rect -206 -181 -149 -180
rect -206 -182 -152 -181
rect -265 -255 -260 -183
rect -206 -184 -205 -182
rect -203 -183 -152 -182
rect -150 -183 -149 -181
rect -127 -182 -121 -180
rect 65 -174 70 -125
rect 96 -123 105 -122
rect 96 -125 98 -123
rect 100 -125 105 -123
rect 96 -126 105 -125
rect 101 -132 105 -126
rect 361 -123 370 -122
rect 361 -125 366 -123
rect 368 -125 370 -123
rect 361 -126 370 -125
rect 396 -123 401 -121
rect 396 -125 398 -123
rect 400 -125 401 -123
rect 504 -123 508 -121
rect 504 -125 505 -123
rect 507 -125 508 -123
rect 139 -132 182 -131
rect 101 -134 179 -132
rect 181 -134 182 -132
rect 101 -135 182 -134
rect 284 -132 327 -131
rect 361 -132 365 -126
rect 284 -134 285 -132
rect 287 -134 365 -132
rect 284 -135 365 -134
rect 101 -137 143 -135
rect 323 -137 365 -135
rect 225 -139 230 -137
rect 225 -141 226 -139
rect 228 -141 230 -139
rect 225 -165 230 -141
rect 225 -167 227 -165
rect 229 -167 230 -165
rect 225 -168 230 -167
rect 236 -139 241 -137
rect 236 -141 238 -139
rect 240 -141 241 -139
rect 236 -165 241 -141
rect 236 -167 238 -165
rect 240 -167 241 -165
rect 236 -168 241 -167
rect 65 -178 71 -174
rect 65 -180 67 -178
rect 69 -180 71 -178
rect 65 -182 71 -180
rect 396 -178 401 -125
rect 405 -126 417 -125
rect 405 -128 406 -126
rect 408 -128 414 -126
rect 416 -128 417 -126
rect 405 -129 417 -128
rect 487 -127 500 -126
rect 487 -129 488 -127
rect 490 -129 495 -127
rect 497 -129 500 -127
rect 487 -130 500 -129
rect 396 -180 398 -178
rect 400 -180 401 -178
rect 396 -181 401 -180
rect -203 -184 -149 -183
rect -206 -185 -149 -184
rect 504 -187 508 -125
rect 534 -123 543 -122
rect 534 -125 536 -123
rect 538 -125 543 -123
rect 534 -126 543 -125
rect 539 -132 543 -126
rect 675 -124 679 -101
rect 691 -115 695 -70
rect 691 -117 692 -115
rect 694 -117 695 -115
rect 691 -118 695 -117
rect 675 -126 676 -124
rect 678 -126 679 -124
rect 699 -123 703 140
rect 823 -9 828 -7
rect 724 -11 828 -9
rect 724 -13 725 -11
rect 727 -13 828 -11
rect 724 -14 828 -13
rect 764 -120 770 -119
rect 699 -125 700 -123
rect 702 -125 703 -123
rect 699 -126 703 -125
rect 756 -123 770 -120
rect 756 -126 757 -123
rect 759 -126 770 -123
rect 675 -129 679 -126
rect 756 -128 770 -126
rect 577 -132 620 -131
rect 539 -134 617 -132
rect 619 -134 620 -132
rect 539 -135 620 -134
rect 539 -137 581 -135
rect 664 -136 672 -134
rect 664 -138 665 -136
rect 667 -138 672 -136
rect 664 -140 672 -138
rect 668 -170 672 -140
rect 668 -173 669 -170
rect 671 -173 672 -170
rect 668 -174 672 -173
rect -72 -189 508 -187
rect -72 -191 -71 -189
rect -69 -191 508 -189
rect -72 -192 508 -191
rect -169 -194 -165 -192
rect -169 -196 -168 -194
rect -166 -196 -165 -194
rect 764 -195 770 -128
rect -169 -224 -165 -196
rect 716 -202 770 -195
rect 588 -211 643 -208
rect 588 -212 638 -211
rect 63 -214 69 -212
rect 63 -216 65 -214
rect 67 -216 69 -214
rect -169 -236 -164 -224
rect 63 -236 69 -216
rect -169 -243 69 -236
rect 418 -213 638 -212
rect 640 -213 643 -211
rect 418 -216 643 -213
rect 418 -217 462 -216
rect 418 -233 423 -217
rect 418 -235 419 -233
rect 421 -235 423 -233
rect 418 -237 423 -235
rect 552 -232 571 -231
rect 552 -233 695 -232
rect 552 -235 554 -233
rect 556 -234 695 -233
rect 556 -235 692 -234
rect 552 -236 692 -235
rect 694 -236 695 -234
rect 552 -237 695 -236
rect 432 -249 595 -245
rect -265 -257 345 -255
rect -265 -259 341 -257
rect 343 -259 345 -257
rect -265 -261 345 -259
rect 432 -257 436 -249
rect 432 -259 433 -257
rect 435 -259 436 -257
rect 432 -260 436 -259
rect 391 -264 404 -263
rect 391 -266 401 -264
rect 403 -266 404 -264
rect 391 -267 404 -266
rect 437 -265 447 -264
rect 437 -267 444 -265
rect 446 -267 447 -265
rect -105 -285 -28 -283
rect -105 -287 -32 -285
rect -30 -287 -28 -285
rect -105 -289 -28 -287
rect -105 -310 -100 -289
rect 391 -303 396 -267
rect 437 -268 447 -267
rect 480 -265 490 -264
rect 480 -267 487 -265
rect 489 -267 490 -265
rect 480 -268 490 -267
rect 437 -294 442 -268
rect 437 -299 473 -294
rect 391 -308 444 -303
rect -105 -312 -104 -310
rect -102 -312 -100 -310
rect -105 -314 -100 -312
rect -261 -341 -248 -340
rect -261 -343 -251 -341
rect -249 -343 -248 -341
rect -261 -344 -248 -343
rect -215 -342 -205 -341
rect -215 -344 -208 -342
rect -206 -344 -205 -342
rect -261 -380 -256 -344
rect -215 -345 -205 -344
rect -172 -342 -162 -341
rect -172 -344 -165 -342
rect -163 -344 -162 -342
rect -172 -345 -162 -344
rect -123 -342 -102 -340
rect -123 -344 -122 -342
rect -120 -344 -102 -342
rect -215 -371 -210 -345
rect -215 -376 -179 -371
rect -261 -385 -208 -380
rect -213 -422 -208 -385
rect -186 -383 -179 -376
rect -172 -373 -167 -345
rect -123 -346 -102 -344
rect -107 -348 -102 -346
rect -83 -346 -29 -340
rect -83 -348 -79 -346
rect -107 -352 -79 -348
rect -107 -353 -102 -352
rect -172 -377 -98 -373
rect -186 -389 -118 -383
rect -213 -424 -212 -422
rect -210 -424 -208 -422
rect -213 -425 -208 -424
rect -126 -430 -120 -389
rect -104 -422 -98 -377
rect -104 -424 -102 -422
rect -100 -424 -98 -422
rect -104 -425 -98 -424
rect -273 -432 -249 -431
rect -126 -432 -124 -430
rect -122 -432 -120 -430
rect -273 -434 -252 -432
rect -250 -434 -249 -432
rect -273 -436 -249 -434
rect -205 -433 -148 -432
rect -205 -434 -151 -433
rect -205 -436 -204 -434
rect -202 -435 -151 -434
rect -149 -435 -148 -433
rect -126 -434 -120 -432
rect -71 -433 -42 -430
rect -202 -436 -148 -435
rect -273 -688 -268 -436
rect -205 -437 -148 -436
rect -71 -435 -70 -433
rect -68 -435 -42 -433
rect -71 -437 -42 -435
rect -168 -445 -164 -443
rect -168 -447 -167 -445
rect -165 -447 -164 -445
rect -168 -481 -164 -447
rect -260 -488 -164 -481
rect -48 -480 -42 -437
rect -48 -482 -46 -480
rect -44 -482 -42 -480
rect -48 -484 -42 -482
rect -260 -676 -255 -488
rect -34 -570 -29 -346
rect 439 -345 444 -308
rect 466 -306 473 -299
rect 480 -296 485 -268
rect 480 -300 554 -296
rect 466 -312 534 -306
rect 439 -347 440 -345
rect 442 -347 444 -345
rect 439 -348 444 -347
rect 526 -353 532 -312
rect 548 -345 554 -300
rect 590 -306 595 -249
rect 590 -308 591 -306
rect 593 -308 595 -306
rect 590 -309 595 -308
rect 548 -347 550 -345
rect 552 -347 554 -345
rect 548 -348 554 -347
rect 388 -354 394 -353
rect 388 -356 403 -354
rect 526 -355 528 -353
rect 530 -355 532 -353
rect 388 -358 400 -356
rect 402 -358 403 -356
rect 388 -360 403 -358
rect 447 -356 504 -355
rect 447 -357 501 -356
rect 447 -359 448 -357
rect 450 -358 501 -357
rect 503 -358 504 -356
rect 526 -357 532 -355
rect 450 -359 504 -358
rect 447 -360 504 -359
rect 388 -408 394 -360
rect 480 -369 496 -367
rect 480 -371 484 -369
rect 486 -371 496 -369
rect 480 -372 496 -371
rect 408 -382 415 -379
rect 408 -384 411 -382
rect 413 -384 415 -382
rect 408 -398 415 -384
rect 408 -400 411 -398
rect 413 -400 415 -398
rect 408 -401 415 -400
rect 491 -394 496 -372
rect 491 -398 500 -394
rect 491 -400 497 -398
rect 499 -400 500 -398
rect 491 -403 500 -400
rect 527 -398 705 -394
rect 527 -400 529 -398
rect 531 -400 705 -398
rect 527 -403 705 -400
rect 388 -410 425 -408
rect 388 -412 422 -410
rect 424 -412 425 -410
rect 388 -414 425 -412
rect 188 -487 331 -482
rect 20 -499 111 -498
rect 147 -499 153 -498
rect 20 -501 21 -499
rect 23 -501 108 -499
rect 110 -501 111 -499
rect 20 -502 111 -501
rect 124 -500 150 -499
rect 124 -502 125 -500
rect 127 -501 150 -500
rect 152 -501 153 -499
rect 127 -502 153 -501
rect 124 -503 153 -502
rect 188 -500 192 -487
rect 188 -502 189 -500
rect 191 -502 192 -500
rect 188 -503 192 -502
rect 286 -492 290 -491
rect 286 -494 287 -492
rect 289 -494 290 -492
rect 286 -500 290 -494
rect 327 -492 331 -487
rect 565 -487 581 -485
rect 565 -489 566 -487
rect 568 -489 581 -487
rect 565 -490 581 -489
rect 327 -494 328 -492
rect 330 -494 331 -492
rect 577 -492 578 -490
rect 580 -492 581 -490
rect 577 -494 581 -492
rect 624 -486 682 -480
rect 327 -495 331 -494
rect 286 -502 287 -500
rect 289 -502 290 -500
rect 286 -503 290 -502
rect 317 -499 323 -498
rect 359 -499 450 -498
rect 317 -501 318 -499
rect 320 -500 346 -499
rect 320 -501 343 -500
rect 317 -502 343 -501
rect 345 -502 346 -500
rect 359 -501 360 -499
rect 362 -501 447 -499
rect 449 -501 450 -499
rect 359 -502 450 -501
rect 458 -499 549 -498
rect 585 -499 591 -498
rect 458 -501 459 -499
rect 461 -501 546 -499
rect 548 -501 549 -499
rect 458 -502 549 -501
rect 562 -500 588 -499
rect 562 -502 563 -500
rect 565 -501 588 -500
rect 590 -501 591 -499
rect 565 -502 591 -501
rect 317 -503 346 -502
rect 562 -503 591 -502
rect 624 -500 629 -486
rect 624 -502 625 -500
rect 627 -502 629 -500
rect 624 -503 629 -502
rect 67 -508 71 -506
rect 67 -510 68 -508
rect 70 -510 71 -508
rect 67 -519 71 -510
rect 98 -508 107 -507
rect 98 -510 100 -508
rect 102 -510 107 -508
rect 98 -511 107 -510
rect 67 -521 68 -519
rect 70 -521 71 -519
rect 67 -522 71 -521
rect 103 -517 107 -511
rect 363 -508 372 -507
rect 363 -510 368 -508
rect 370 -510 372 -508
rect 363 -511 372 -510
rect 399 -508 403 -507
rect 399 -510 400 -508
rect 402 -510 403 -508
rect 141 -517 184 -516
rect 103 -519 181 -517
rect 183 -519 184 -517
rect 103 -520 184 -519
rect 286 -517 329 -516
rect 363 -517 367 -511
rect 286 -519 287 -517
rect 289 -519 367 -517
rect 286 -520 367 -519
rect 103 -522 145 -520
rect 325 -522 367 -520
rect 399 -519 403 -510
rect 505 -508 509 -506
rect 505 -510 506 -508
rect 508 -510 509 -508
rect 399 -521 400 -519
rect 402 -521 403 -519
rect 409 -515 414 -511
rect 409 -516 419 -515
rect 409 -518 410 -516
rect 412 -518 416 -516
rect 418 -518 419 -516
rect 409 -520 419 -518
rect 489 -517 500 -516
rect 489 -519 490 -517
rect 492 -519 497 -517
rect 499 -519 500 -517
rect 489 -520 500 -519
rect 399 -522 403 -521
rect 505 -521 509 -510
rect 536 -508 545 -507
rect 536 -510 538 -508
rect 540 -510 545 -508
rect 536 -511 545 -510
rect 227 -524 232 -522
rect 227 -526 228 -524
rect 230 -526 232 -524
rect -34 -571 188 -570
rect -34 -573 184 -571
rect 186 -573 188 -571
rect -34 -575 188 -573
rect 227 -571 232 -526
rect 227 -573 229 -571
rect 231 -573 232 -571
rect 227 -576 232 -573
rect 238 -524 243 -522
rect 238 -526 240 -524
rect 242 -526 243 -524
rect 505 -523 506 -521
rect 508 -523 509 -521
rect 541 -517 545 -511
rect 677 -509 681 -486
rect 677 -511 678 -509
rect 680 -511 681 -509
rect 701 -508 705 -403
rect 717 -500 722 -202
rect 823 -208 828 -14
rect 772 -211 828 -208
rect 772 -213 775 -211
rect 777 -213 828 -211
rect 772 -216 828 -213
rect 823 -217 828 -216
rect 717 -502 718 -500
rect 720 -502 722 -500
rect 717 -503 722 -502
rect 701 -510 702 -508
rect 704 -510 705 -508
rect 701 -511 705 -510
rect 677 -514 681 -511
rect 579 -517 622 -516
rect 541 -519 619 -517
rect 621 -519 622 -517
rect 541 -520 622 -519
rect 541 -522 583 -520
rect 505 -526 509 -523
rect 238 -571 243 -526
rect 452 -559 456 -557
rect 452 -561 453 -559
rect 455 -561 456 -559
rect 238 -576 448 -571
rect -79 -621 64 -616
rect -247 -633 -156 -632
rect -120 -633 -114 -632
rect -247 -635 -246 -633
rect -244 -635 -159 -633
rect -157 -635 -156 -633
rect -247 -636 -156 -635
rect -143 -634 -117 -633
rect -143 -636 -142 -634
rect -140 -635 -117 -634
rect -115 -635 -114 -633
rect -140 -636 -114 -635
rect -143 -637 -114 -636
rect -79 -634 -75 -621
rect -79 -636 -78 -634
rect -76 -636 -75 -634
rect -79 -637 -75 -636
rect 19 -626 23 -625
rect 19 -628 20 -626
rect 22 -628 23 -626
rect 19 -634 23 -628
rect 60 -626 64 -621
rect 298 -621 314 -619
rect 298 -623 299 -621
rect 301 -623 314 -621
rect 298 -624 314 -623
rect 60 -628 61 -626
rect 63 -628 64 -626
rect 310 -626 311 -624
rect 313 -626 314 -624
rect 310 -628 314 -626
rect 357 -620 415 -614
rect 60 -629 64 -628
rect 19 -636 20 -634
rect 22 -636 23 -634
rect 19 -637 23 -636
rect 50 -633 56 -632
rect 92 -633 183 -632
rect 50 -635 51 -633
rect 53 -634 79 -633
rect 53 -635 76 -634
rect 50 -636 76 -635
rect 78 -636 79 -634
rect 92 -635 93 -633
rect 95 -635 180 -633
rect 182 -635 183 -633
rect 92 -636 183 -635
rect 191 -633 282 -632
rect 318 -633 324 -632
rect 191 -635 192 -633
rect 194 -635 279 -633
rect 281 -635 282 -633
rect 191 -636 282 -635
rect 295 -634 321 -633
rect 295 -636 296 -634
rect 298 -635 321 -634
rect 323 -635 324 -633
rect 298 -636 324 -635
rect 50 -637 79 -636
rect 295 -637 324 -636
rect 357 -634 362 -620
rect 357 -636 358 -634
rect 360 -636 362 -634
rect 357 -637 362 -636
rect -200 -642 -196 -640
rect -200 -644 -199 -642
rect -197 -644 -196 -642
rect -223 -651 -212 -650
rect -223 -653 -222 -651
rect -220 -653 -215 -651
rect -213 -653 -212 -651
rect -223 -654 -212 -653
rect -200 -676 -196 -644
rect -169 -642 -160 -641
rect -169 -644 -167 -642
rect -165 -644 -160 -642
rect -169 -645 -160 -644
rect -164 -651 -160 -645
rect 96 -642 105 -641
rect 96 -644 101 -642
rect 103 -644 105 -642
rect 96 -645 105 -644
rect 127 -642 132 -640
rect 127 -644 129 -642
rect 131 -644 132 -642
rect -126 -651 -83 -650
rect -164 -653 -86 -651
rect -84 -653 -83 -651
rect -164 -654 -83 -653
rect 19 -651 62 -650
rect 96 -651 100 -645
rect 19 -653 20 -651
rect 22 -653 100 -651
rect 19 -654 100 -653
rect -164 -656 -122 -654
rect 58 -656 100 -654
rect -260 -683 -196 -676
rect 127 -688 132 -644
rect 239 -642 243 -640
rect 239 -644 240 -642
rect 242 -644 243 -642
rect 216 -646 220 -645
rect 216 -648 217 -646
rect 219 -648 220 -646
rect 216 -649 220 -648
rect 148 -651 152 -649
rect 148 -653 149 -651
rect 151 -653 152 -651
rect 148 -669 152 -653
rect 216 -651 226 -649
rect 216 -653 223 -651
rect 225 -653 226 -651
rect 216 -654 226 -653
rect 216 -655 220 -654
rect 148 -671 149 -669
rect 151 -671 152 -669
rect 148 -672 152 -671
rect -273 -696 132 -688
rect 239 -680 243 -644
rect 269 -642 278 -641
rect 269 -644 271 -642
rect 273 -644 278 -642
rect 269 -645 278 -644
rect 274 -651 278 -645
rect 410 -643 414 -620
rect 410 -645 411 -643
rect 413 -645 414 -643
rect 444 -642 448 -576
rect 452 -634 456 -561
rect 452 -636 453 -634
rect 455 -636 456 -634
rect 452 -637 456 -636
rect 444 -644 445 -642
rect 447 -644 448 -642
rect 444 -645 448 -644
rect 410 -648 414 -645
rect 312 -651 355 -650
rect 274 -653 352 -651
rect 354 -653 355 -651
rect 274 -654 355 -653
rect 274 -656 316 -654
rect 239 -707 244 -680
rect 4 -708 244 -707
rect 4 -710 5 -708
rect 7 -710 244 -708
rect 4 -712 244 -710
<< alu3 >>
rect -33 199 -28 201
rect -33 197 -31 199
rect -29 197 -28 199
rect -33 -285 -28 197
rect 493 55 500 57
rect 493 53 495 55
rect 497 53 500 55
rect 251 7 393 8
rect 251 5 253 7
rect 255 6 393 7
rect 255 5 388 6
rect 251 4 388 5
rect 391 4 393 6
rect 251 3 393 4
rect 55 -9 355 -8
rect 55 -11 352 -9
rect 354 -11 355 -9
rect 55 -13 355 -11
rect 55 -15 60 -13
rect 55 -132 59 -15
rect 493 -38 500 53
rect 687 -10 728 -9
rect 687 -12 688 -10
rect 690 -11 728 -10
rect 690 -12 725 -11
rect 687 -13 725 -12
rect 727 -13 728 -11
rect 687 -14 728 -13
rect 651 -27 816 -23
rect 651 -29 654 -27
rect 656 -29 816 -27
rect 651 -32 816 -29
rect 493 -40 495 -38
rect 497 -40 500 -38
rect 493 -42 500 -40
rect 55 -134 56 -132
rect 58 -134 59 -132
rect 55 -135 59 -134
rect 140 -99 144 -98
rect 140 -101 141 -99
rect 143 -101 144 -99
rect 65 -177 71 -174
rect 63 -178 71 -177
rect 63 -180 67 -178
rect 69 -180 71 -178
rect 63 -184 71 -180
rect 63 -214 69 -184
rect 63 -216 65 -214
rect 67 -216 69 -214
rect 63 -218 69 -216
rect -33 -287 -32 -285
rect -30 -287 -28 -285
rect -33 -289 -28 -287
rect -1 -369 4 -368
rect 140 -369 144 -101
rect 555 -102 567 -100
rect 555 -104 564 -102
rect 566 -104 567 -102
rect 555 -105 567 -104
rect 284 -107 559 -105
rect 284 -109 285 -107
rect 287 -109 559 -107
rect 284 -110 559 -109
rect 405 -115 410 -114
rect 405 -117 406 -115
rect 408 -117 410 -115
rect 405 -126 410 -117
rect 405 -128 406 -126
rect 408 -128 410 -126
rect 405 -129 410 -128
rect 492 -115 500 -114
rect 492 -117 495 -115
rect 497 -117 500 -115
rect 492 -127 500 -117
rect 492 -129 495 -127
rect 497 -129 500 -127
rect 492 -130 500 -129
rect -1 -376 144 -369
rect 225 -165 230 -163
rect 225 -167 227 -165
rect 229 -167 230 -165
rect -1 -377 141 -376
rect -48 -480 -42 -477
rect -48 -482 -46 -480
rect -44 -482 -42 -480
rect -48 -524 -42 -482
rect -48 -526 -47 -524
rect -45 -526 -42 -524
rect -48 -530 -42 -526
rect -1 -584 4 -377
rect 225 -408 230 -167
rect 59 -414 230 -408
rect 236 -165 241 -163
rect 236 -167 238 -165
rect 240 -167 241 -165
rect 236 -408 241 -167
rect 668 -170 672 -168
rect 668 -173 669 -170
rect 671 -173 672 -170
rect 391 -178 401 -176
rect 391 -180 398 -178
rect 400 -180 401 -178
rect 391 -181 401 -180
rect 391 -203 396 -181
rect 340 -209 396 -203
rect 340 -257 345 -209
rect 340 -259 341 -257
rect 343 -259 345 -257
rect 340 -261 345 -259
rect 408 -398 415 -396
rect 408 -400 411 -398
rect 413 -400 415 -398
rect 236 -410 388 -408
rect 236 -412 385 -410
rect 387 -412 388 -410
rect 236 -414 388 -412
rect 59 -518 63 -414
rect 408 -456 415 -400
rect 496 -398 500 -394
rect 496 -400 497 -398
rect 499 -400 500 -398
rect 420 -410 492 -408
rect 420 -412 422 -410
rect 424 -412 492 -410
rect 420 -414 492 -412
rect 487 -426 492 -414
rect 496 -416 500 -400
rect 496 -418 497 -416
rect 499 -418 500 -416
rect 496 -420 500 -418
rect 528 -398 532 -394
rect 528 -400 529 -398
rect 531 -400 532 -398
rect 528 -426 532 -400
rect 487 -430 532 -426
rect 514 -448 528 -447
rect 668 -448 672 -173
rect 691 -234 695 -232
rect 691 -236 692 -234
rect 694 -236 695 -234
rect 691 -256 695 -236
rect 809 -255 816 -32
rect 708 -256 816 -255
rect 691 -266 816 -256
rect 809 -267 816 -266
rect 514 -449 672 -448
rect 514 -451 516 -449
rect 518 -451 672 -449
rect 514 -453 672 -451
rect 408 -458 410 -456
rect 412 -458 415 -456
rect 408 -461 415 -458
rect 557 -487 569 -485
rect 557 -489 566 -487
rect 568 -489 569 -487
rect 557 -490 569 -489
rect 286 -492 561 -490
rect 286 -494 287 -492
rect 289 -494 561 -492
rect 286 -495 561 -494
rect 409 -502 414 -500
rect 409 -504 410 -502
rect 412 -504 414 -502
rect 409 -516 414 -504
rect 409 -518 410 -516
rect 412 -518 414 -516
rect 59 -519 71 -518
rect 59 -521 68 -519
rect 70 -521 71 -519
rect 59 -522 71 -521
rect 383 -519 403 -518
rect 383 -521 384 -519
rect 386 -521 400 -519
rect 402 -521 403 -519
rect 409 -520 414 -518
rect 496 -506 500 -505
rect 496 -508 497 -506
rect 499 -508 500 -506
rect 496 -517 500 -508
rect 496 -519 497 -517
rect 499 -519 500 -517
rect 496 -520 500 -519
rect 383 -522 403 -521
rect 505 -521 519 -520
rect 505 -523 506 -521
rect 508 -522 519 -521
rect 508 -523 515 -522
rect 505 -524 515 -523
rect 517 -524 519 -522
rect 505 -526 519 -524
rect 182 -559 456 -557
rect 182 -561 453 -559
rect 455 -561 456 -559
rect 182 -562 456 -561
rect 182 -571 188 -562
rect 182 -573 184 -571
rect 186 -573 188 -571
rect 182 -575 188 -573
rect 227 -571 232 -568
rect 227 -573 229 -571
rect 231 -573 232 -571
rect -223 -589 4 -584
rect 227 -588 232 -573
rect -223 -651 -219 -589
rect 227 -590 228 -588
rect 230 -590 232 -588
rect 227 -592 232 -590
rect 290 -621 302 -619
rect 290 -623 299 -621
rect 301 -623 302 -621
rect 290 -624 302 -623
rect 19 -626 294 -624
rect 19 -628 20 -626
rect 22 -628 294 -626
rect 19 -629 294 -628
rect 216 -637 220 -635
rect 216 -639 217 -637
rect 219 -639 220 -637
rect 216 -646 220 -639
rect 216 -648 217 -646
rect 219 -648 220 -646
rect 216 -649 220 -648
rect -223 -653 -222 -651
rect -220 -653 -219 -651
rect -223 -654 -219 -653
rect -48 -708 9 -705
rect -48 -710 -47 -708
rect -45 -710 5 -708
rect 7 -710 9 -708
rect -48 -712 9 -710
<< alu4 >>
rect 386 6 393 8
rect 386 4 388 6
rect 391 4 393 6
rect 386 -113 393 4
rect 493 -38 500 -36
rect 493 -40 495 -38
rect 497 -40 500 -38
rect 386 -115 411 -113
rect 386 -117 406 -115
rect 408 -117 411 -115
rect 386 -120 411 -117
rect 493 -115 500 -40
rect 493 -117 495 -115
rect 497 -117 500 -115
rect 493 -118 500 -117
rect 383 -410 389 -408
rect 383 -412 385 -410
rect 387 -412 389 -410
rect 383 -519 389 -412
rect 496 -416 500 -414
rect 496 -418 497 -416
rect 499 -418 500 -416
rect 408 -456 415 -453
rect 408 -458 410 -456
rect 412 -458 415 -456
rect 408 -461 415 -458
rect 409 -502 414 -461
rect 409 -504 410 -502
rect 412 -504 414 -502
rect 409 -506 414 -504
rect 496 -506 500 -418
rect 496 -508 497 -506
rect 499 -508 500 -506
rect 496 -510 500 -508
rect 514 -449 519 -447
rect 514 -451 516 -449
rect 518 -451 519 -449
rect 383 -521 384 -519
rect 386 -521 389 -519
rect -48 -524 -44 -521
rect 383 -522 389 -521
rect 514 -522 519 -451
rect -48 -526 -47 -524
rect -45 -526 -44 -524
rect 514 -524 515 -522
rect 517 -524 519 -522
rect 514 -526 519 -524
rect -48 -708 -44 -526
rect 227 -586 232 -584
rect 216 -588 232 -586
rect 216 -590 228 -588
rect 230 -590 232 -588
rect 216 -592 232 -590
rect 216 -597 221 -592
rect 216 -637 220 -597
rect 216 -639 217 -637
rect 219 -639 220 -637
rect 216 -640 220 -639
rect -48 -710 -47 -708
rect -45 -710 -44 -708
rect -48 -712 -44 -710
<< ptie >>
rect -252 -108 -246 -106
rect -252 -110 -250 -108
rect -248 -110 -246 -108
rect -252 -112 -246 -110
rect -209 -108 -203 -106
rect -209 -110 -207 -108
rect -205 -110 -203 -108
rect -209 -112 -203 -110
rect -166 -108 -160 -106
rect -166 -110 -164 -108
rect -162 -110 -160 -108
rect -166 -112 -160 -110
rect -123 -108 -117 -106
rect -123 -110 -121 -108
rect -119 -110 -117 -108
rect -123 -112 -117 -110
rect -251 -360 -245 -358
rect -251 -362 -249 -360
rect -247 -362 -245 -360
rect -251 -364 -245 -362
rect -208 -360 -202 -358
rect -208 -362 -206 -360
rect -204 -362 -202 -360
rect -208 -364 -202 -362
rect -165 -360 -159 -358
rect -165 -362 -163 -360
rect -161 -362 -159 -360
rect -165 -364 -159 -362
rect -122 -360 -116 -358
rect -122 -362 -120 -360
rect -118 -362 -116 -360
rect -122 -364 -116 -362
rect 268 134 274 136
rect 268 132 270 134
rect 272 132 274 134
rect 268 130 274 132
rect 311 134 317 136
rect 311 132 313 134
rect 315 132 317 134
rect 311 130 317 132
rect 354 134 360 136
rect 354 132 356 134
rect 358 132 360 134
rect 354 130 360 132
rect 397 134 403 136
rect 397 132 399 134
rect 401 132 403 134
rect 397 130 403 132
rect 106 -149 140 -147
rect 106 -151 108 -149
rect 110 -151 136 -149
rect 138 -151 140 -149
rect 106 -153 140 -151
rect 326 -149 360 -147
rect 326 -151 328 -149
rect 330 -151 356 -149
rect 358 -151 360 -149
rect 326 -153 360 -151
rect 544 -149 578 -147
rect 544 -151 546 -149
rect 548 -151 574 -149
rect 576 -151 578 -149
rect 544 -153 578 -151
rect 401 -283 407 -281
rect 401 -285 403 -283
rect 405 -285 407 -283
rect 401 -287 407 -285
rect 444 -283 450 -281
rect 444 -285 446 -283
rect 448 -285 450 -283
rect 444 -287 450 -285
rect 487 -283 493 -281
rect 487 -285 489 -283
rect 491 -285 493 -283
rect 487 -287 493 -285
rect 530 -283 536 -281
rect 530 -285 532 -283
rect 534 -285 536 -283
rect 530 -287 536 -285
rect 108 -534 142 -532
rect 108 -536 110 -534
rect 112 -536 138 -534
rect 140 -536 142 -534
rect 108 -538 142 -536
rect 328 -534 362 -532
rect 328 -536 330 -534
rect 332 -536 358 -534
rect 360 -536 362 -534
rect 328 -538 362 -536
rect 546 -534 580 -532
rect 546 -536 548 -534
rect 550 -536 576 -534
rect 578 -536 580 -534
rect 546 -538 580 -536
rect -159 -668 -125 -666
rect -159 -670 -157 -668
rect -155 -670 -129 -668
rect -127 -670 -125 -668
rect -159 -672 -125 -670
rect 61 -668 95 -666
rect 61 -670 63 -668
rect 65 -670 91 -668
rect 93 -670 95 -668
rect 61 -672 95 -670
rect 279 -668 313 -666
rect 279 -670 281 -668
rect 283 -670 309 -668
rect 311 -670 313 -668
rect 279 -672 313 -670
<< ntie >>
rect 268 194 302 196
rect 268 192 270 194
rect 272 192 284 194
rect 286 192 298 194
rect 300 192 302 194
rect 268 190 302 192
rect 311 194 345 196
rect 311 192 313 194
rect 315 192 327 194
rect 329 192 341 194
rect 343 192 345 194
rect 311 190 345 192
rect 354 194 388 196
rect 354 192 356 194
rect 358 192 370 194
rect 372 192 384 194
rect 386 192 388 194
rect 354 190 388 192
rect 397 194 431 196
rect 397 192 399 194
rect 401 192 413 194
rect 415 192 427 194
rect 429 192 431 194
rect 397 190 431 192
rect -252 -48 -218 -46
rect -252 -50 -250 -48
rect -248 -50 -236 -48
rect -234 -50 -222 -48
rect -220 -50 -218 -48
rect -252 -52 -218 -50
rect -209 -48 -175 -46
rect -209 -50 -207 -48
rect -205 -50 -193 -48
rect -191 -50 -179 -48
rect -177 -50 -175 -48
rect -209 -52 -175 -50
rect -166 -48 -132 -46
rect -166 -50 -164 -48
rect -162 -50 -150 -48
rect -148 -50 -136 -48
rect -134 -50 -132 -48
rect -166 -52 -132 -50
rect -123 -48 -89 -46
rect -123 -50 -121 -48
rect -119 -50 -107 -48
rect -105 -50 -93 -48
rect -91 -50 -89 -48
rect -123 -52 -89 -50
rect -251 -300 -217 -298
rect -251 -302 -249 -300
rect -247 -302 -235 -300
rect -233 -302 -221 -300
rect -219 -302 -217 -300
rect -251 -304 -217 -302
rect -208 -300 -174 -298
rect -208 -302 -206 -300
rect -204 -302 -192 -300
rect -190 -302 -178 -300
rect -176 -302 -174 -300
rect -208 -304 -174 -302
rect -165 -300 -131 -298
rect -165 -302 -163 -300
rect -161 -302 -149 -300
rect -147 -302 -135 -300
rect -133 -302 -131 -300
rect -165 -304 -131 -302
rect -122 -300 -88 -298
rect -122 -302 -120 -300
rect -118 -302 -106 -300
rect -104 -302 -92 -300
rect -90 -302 -88 -300
rect -122 -304 -88 -302
rect 134 -89 140 -87
rect 134 -91 136 -89
rect 138 -91 140 -89
rect 134 -93 140 -91
rect 326 -89 332 -87
rect 326 -91 328 -89
rect 330 -91 332 -89
rect 326 -93 332 -91
rect 572 -89 578 -87
rect 572 -91 574 -89
rect 576 -91 578 -89
rect 572 -93 578 -91
rect 401 -223 435 -221
rect 401 -225 403 -223
rect 405 -225 417 -223
rect 419 -225 431 -223
rect 433 -225 435 -223
rect 401 -227 435 -225
rect 444 -223 478 -221
rect 444 -225 446 -223
rect 448 -225 460 -223
rect 462 -225 474 -223
rect 476 -225 478 -223
rect 444 -227 478 -225
rect 487 -223 521 -221
rect 487 -225 489 -223
rect 491 -225 503 -223
rect 505 -225 517 -223
rect 519 -225 521 -223
rect 487 -227 521 -225
rect 530 -223 564 -221
rect 530 -225 532 -223
rect 534 -225 546 -223
rect 548 -225 560 -223
rect 562 -225 564 -223
rect 530 -227 564 -225
rect 136 -474 142 -472
rect 136 -476 138 -474
rect 140 -476 142 -474
rect 136 -478 142 -476
rect 328 -474 334 -472
rect 328 -476 330 -474
rect 332 -476 334 -474
rect 328 -478 334 -476
rect 574 -474 580 -472
rect 574 -476 576 -474
rect 578 -476 580 -474
rect 574 -478 580 -476
rect -131 -608 -125 -606
rect -131 -610 -129 -608
rect -127 -610 -125 -608
rect -131 -612 -125 -610
rect 61 -608 67 -606
rect 61 -610 63 -608
rect 65 -610 67 -608
rect 61 -612 67 -610
rect 307 -608 313 -606
rect 307 -610 309 -608
rect 311 -610 313 -608
rect 307 -612 313 -610
<< nmos >>
rect -246 -100 -244 -94
rect -234 -106 -232 -97
rect -227 -106 -225 -97
rect -203 -100 -201 -94
rect -191 -106 -189 -97
rect -184 -106 -182 -97
rect -160 -100 -158 -94
rect -148 -106 -146 -97
rect -141 -106 -139 -97
rect -117 -100 -115 -94
rect -105 -106 -103 -97
rect -98 -106 -96 -97
rect -247 -205 -245 -192
rect -237 -202 -235 -192
rect -227 -199 -225 -185
rect -217 -199 -215 -185
rect -197 -205 -195 -185
rect -190 -205 -188 -185
rect -179 -205 -177 -191
rect -145 -205 -143 -191
rect -134 -205 -132 -185
rect -127 -205 -125 -185
rect -107 -199 -105 -185
rect -97 -199 -95 -185
rect -87 -202 -85 -192
rect -77 -205 -75 -192
rect -245 -352 -243 -346
rect -233 -358 -231 -349
rect -226 -358 -224 -349
rect -202 -352 -200 -346
rect -190 -358 -188 -349
rect -183 -358 -181 -349
rect -159 -352 -157 -346
rect -147 -358 -145 -349
rect -140 -358 -138 -349
rect -116 -352 -114 -346
rect -104 -358 -102 -349
rect -97 -358 -95 -349
rect 274 142 276 148
rect 286 136 288 145
rect 293 136 295 145
rect 317 142 319 148
rect 329 136 331 145
rect 336 136 338 145
rect 360 142 362 148
rect 372 136 374 145
rect 379 136 381 145
rect 403 142 405 148
rect 415 136 417 145
rect 422 136 424 145
rect 273 37 275 50
rect 283 40 285 50
rect 293 43 295 57
rect 303 43 305 57
rect 323 37 325 57
rect 330 37 332 57
rect 341 37 343 51
rect 375 37 377 51
rect 386 37 388 57
rect 393 37 395 57
rect 413 43 415 57
rect 423 43 425 57
rect 433 40 435 50
rect 443 37 445 50
rect 24 -150 26 -136
rect 35 -150 37 -130
rect 42 -150 44 -130
rect 62 -144 64 -130
rect 72 -144 74 -130
rect 82 -147 84 -137
rect 92 -150 94 -137
rect 112 -141 114 -135
rect 122 -141 124 -135
rect 132 -141 134 -135
rect 153 -150 155 -136
rect 164 -150 166 -130
rect 171 -150 173 -130
rect 191 -144 193 -130
rect 201 -144 203 -130
rect 211 -147 213 -137
rect 221 -150 223 -137
rect 243 -150 245 -137
rect 253 -147 255 -137
rect 263 -144 265 -130
rect 273 -144 275 -130
rect 293 -150 295 -130
rect 300 -150 302 -130
rect 311 -150 313 -136
rect 332 -141 334 -135
rect 342 -141 344 -135
rect 352 -141 354 -135
rect 372 -150 374 -137
rect 382 -147 384 -137
rect 392 -144 394 -130
rect 402 -144 404 -130
rect 422 -150 424 -130
rect 429 -150 431 -130
rect 440 -150 442 -136
rect 462 -150 464 -136
rect 473 -150 475 -130
rect 480 -150 482 -130
rect 500 -144 502 -130
rect 510 -144 512 -130
rect 520 -147 522 -137
rect 530 -150 532 -137
rect 550 -141 552 -135
rect 560 -141 562 -135
rect 570 -141 572 -135
rect 591 -150 593 -136
rect 602 -150 604 -130
rect 609 -150 611 -130
rect 629 -144 631 -130
rect 639 -144 641 -130
rect 649 -147 651 -137
rect 659 -150 661 -137
rect 683 -150 685 -136
rect 694 -150 696 -130
rect 701 -150 703 -130
rect 721 -144 723 -130
rect 731 -144 733 -130
rect 741 -147 743 -137
rect 751 -150 753 -137
rect 407 -275 409 -269
rect 419 -281 421 -272
rect 426 -281 428 -272
rect 450 -275 452 -269
rect 462 -281 464 -272
rect 469 -281 471 -272
rect 493 -275 495 -269
rect 505 -281 507 -272
rect 512 -281 514 -272
rect 536 -275 538 -269
rect 548 -281 550 -272
rect 555 -281 557 -272
rect 406 -380 408 -367
rect 416 -377 418 -367
rect 426 -374 428 -360
rect 436 -374 438 -360
rect 456 -380 458 -360
rect 463 -380 465 -360
rect 474 -380 476 -366
rect 508 -380 510 -366
rect 519 -380 521 -360
rect 526 -380 528 -360
rect 546 -374 548 -360
rect 556 -374 558 -360
rect 566 -377 568 -367
rect 576 -380 578 -367
rect -246 -457 -244 -444
rect -236 -454 -234 -444
rect -226 -451 -224 -437
rect -216 -451 -214 -437
rect -196 -457 -194 -437
rect -189 -457 -187 -437
rect -178 -457 -176 -443
rect -144 -457 -142 -443
rect -133 -457 -131 -437
rect -126 -457 -124 -437
rect -106 -451 -104 -437
rect -96 -451 -94 -437
rect -86 -454 -84 -444
rect -76 -457 -74 -444
rect 26 -535 28 -521
rect 37 -535 39 -515
rect 44 -535 46 -515
rect 64 -529 66 -515
rect 74 -529 76 -515
rect 84 -532 86 -522
rect 94 -535 96 -522
rect 114 -526 116 -520
rect 124 -526 126 -520
rect 134 -526 136 -520
rect 155 -535 157 -521
rect 166 -535 168 -515
rect 173 -535 175 -515
rect 193 -529 195 -515
rect 203 -529 205 -515
rect 213 -532 215 -522
rect 223 -535 225 -522
rect 245 -535 247 -522
rect 255 -532 257 -522
rect 265 -529 267 -515
rect 275 -529 277 -515
rect 295 -535 297 -515
rect 302 -535 304 -515
rect 313 -535 315 -521
rect 334 -526 336 -520
rect 344 -526 346 -520
rect 354 -526 356 -520
rect 374 -535 376 -522
rect 384 -532 386 -522
rect 394 -529 396 -515
rect 404 -529 406 -515
rect 424 -535 426 -515
rect 431 -535 433 -515
rect 442 -535 444 -521
rect 464 -535 466 -521
rect 475 -535 477 -515
rect 482 -535 484 -515
rect 502 -529 504 -515
rect 512 -529 514 -515
rect 522 -532 524 -522
rect 532 -535 534 -522
rect 552 -526 554 -520
rect 562 -526 564 -520
rect 572 -526 574 -520
rect 593 -535 595 -521
rect 604 -535 606 -515
rect 611 -535 613 -515
rect 631 -529 633 -515
rect 641 -529 643 -515
rect 651 -532 653 -522
rect 661 -535 663 -522
rect 685 -535 687 -521
rect 696 -535 698 -515
rect 703 -535 705 -515
rect 723 -529 725 -515
rect 733 -529 735 -515
rect 743 -532 745 -522
rect 753 -535 755 -522
rect -241 -669 -239 -655
rect -230 -669 -228 -649
rect -223 -669 -221 -649
rect -203 -663 -201 -649
rect -193 -663 -191 -649
rect -183 -666 -181 -656
rect -173 -669 -171 -656
rect -153 -660 -151 -654
rect -143 -660 -141 -654
rect -133 -660 -131 -654
rect -112 -669 -110 -655
rect -101 -669 -99 -649
rect -94 -669 -92 -649
rect -74 -663 -72 -649
rect -64 -663 -62 -649
rect -54 -666 -52 -656
rect -44 -669 -42 -656
rect -22 -669 -20 -656
rect -12 -666 -10 -656
rect -2 -663 0 -649
rect 8 -663 10 -649
rect 28 -669 30 -649
rect 35 -669 37 -649
rect 46 -669 48 -655
rect 67 -660 69 -654
rect 77 -660 79 -654
rect 87 -660 89 -654
rect 107 -669 109 -656
rect 117 -666 119 -656
rect 127 -663 129 -649
rect 137 -663 139 -649
rect 157 -669 159 -649
rect 164 -669 166 -649
rect 175 -669 177 -655
rect 197 -669 199 -655
rect 208 -669 210 -649
rect 215 -669 217 -649
rect 235 -663 237 -649
rect 245 -663 247 -649
rect 255 -666 257 -656
rect 265 -669 267 -656
rect 285 -660 287 -654
rect 295 -660 297 -654
rect 305 -660 307 -654
rect 326 -669 328 -655
rect 337 -669 339 -649
rect 344 -669 346 -649
rect 364 -663 366 -649
rect 374 -663 376 -649
rect 384 -666 386 -656
rect 394 -669 396 -656
rect 418 -669 420 -655
rect 429 -669 431 -649
rect 436 -669 438 -649
rect 456 -663 458 -649
rect 466 -663 468 -649
rect 476 -666 478 -656
rect 486 -669 488 -656
<< pmos >>
rect -246 -77 -244 -65
rect -236 -77 -234 -67
rect -226 -77 -224 -67
rect -203 -77 -201 -65
rect -193 -77 -191 -67
rect -183 -77 -181 -67
rect -160 -77 -158 -65
rect -150 -77 -148 -67
rect -140 -77 -138 -67
rect -117 -77 -115 -65
rect -107 -77 -105 -67
rect -97 -77 -95 -67
rect -247 -170 -245 -145
rect -234 -170 -232 -157
rect -224 -173 -222 -148
rect -217 -173 -215 -148
rect -199 -173 -197 -145
rect -189 -173 -187 -145
rect -179 -173 -177 -145
rect -145 -173 -143 -145
rect -135 -173 -133 -145
rect -125 -173 -123 -145
rect -107 -173 -105 -148
rect -100 -173 -98 -148
rect -90 -170 -88 -157
rect -77 -170 -75 -145
rect -245 -329 -243 -317
rect -235 -329 -233 -319
rect -225 -329 -223 -319
rect -202 -329 -200 -317
rect -192 -329 -190 -319
rect -182 -329 -180 -319
rect -159 -329 -157 -317
rect -149 -329 -147 -319
rect -139 -329 -137 -319
rect -116 -329 -114 -317
rect -106 -329 -104 -319
rect -96 -329 -94 -319
rect 274 165 276 177
rect 284 165 286 175
rect 294 165 296 175
rect 317 165 319 177
rect 327 165 329 175
rect 337 165 339 175
rect 360 165 362 177
rect 370 165 372 175
rect 380 165 382 175
rect 403 165 405 177
rect 413 165 415 175
rect 423 165 425 175
rect 273 72 275 97
rect 286 72 288 85
rect 296 69 298 94
rect 303 69 305 94
rect 321 69 323 97
rect 331 69 333 97
rect 341 69 343 97
rect 375 69 377 97
rect 385 69 387 97
rect 395 69 397 97
rect 413 69 415 94
rect 420 69 422 94
rect 430 72 432 85
rect 443 72 445 97
rect 24 -118 26 -90
rect 34 -118 36 -90
rect 44 -118 46 -90
rect 62 -118 64 -93
rect 69 -118 71 -93
rect 79 -115 81 -102
rect 92 -115 94 -90
rect 112 -108 114 -90
rect 119 -108 121 -90
rect 132 -111 134 -99
rect 153 -118 155 -90
rect 163 -118 165 -90
rect 173 -118 175 -90
rect 191 -118 193 -93
rect 198 -118 200 -93
rect 208 -115 210 -102
rect 221 -115 223 -90
rect 243 -115 245 -90
rect 256 -115 258 -102
rect 266 -118 268 -93
rect 273 -118 275 -93
rect 291 -118 293 -90
rect 301 -118 303 -90
rect 311 -118 313 -90
rect 332 -111 334 -99
rect 345 -108 347 -90
rect 352 -108 354 -90
rect 372 -115 374 -90
rect 385 -115 387 -102
rect 395 -118 397 -93
rect 402 -118 404 -93
rect 420 -118 422 -90
rect 430 -118 432 -90
rect 440 -118 442 -90
rect 462 -118 464 -90
rect 472 -118 474 -90
rect 482 -118 484 -90
rect 500 -118 502 -93
rect 507 -118 509 -93
rect 517 -115 519 -102
rect 530 -115 532 -90
rect 550 -108 552 -90
rect 557 -108 559 -90
rect 570 -111 572 -99
rect 591 -118 593 -90
rect 601 -118 603 -90
rect 611 -118 613 -90
rect 629 -118 631 -93
rect 636 -118 638 -93
rect 646 -115 648 -102
rect 659 -115 661 -90
rect 683 -118 685 -90
rect 693 -118 695 -90
rect 703 -118 705 -90
rect 721 -118 723 -93
rect 728 -118 730 -93
rect 738 -115 740 -102
rect 751 -115 753 -90
rect 407 -252 409 -240
rect 417 -252 419 -242
rect 427 -252 429 -242
rect 450 -252 452 -240
rect 460 -252 462 -242
rect 470 -252 472 -242
rect 493 -252 495 -240
rect 503 -252 505 -242
rect 513 -252 515 -242
rect 536 -252 538 -240
rect 546 -252 548 -242
rect 556 -252 558 -242
rect 406 -345 408 -320
rect 419 -345 421 -332
rect 429 -348 431 -323
rect 436 -348 438 -323
rect 454 -348 456 -320
rect 464 -348 466 -320
rect 474 -348 476 -320
rect 508 -348 510 -320
rect 518 -348 520 -320
rect 528 -348 530 -320
rect 546 -348 548 -323
rect 553 -348 555 -323
rect 563 -345 565 -332
rect 576 -345 578 -320
rect -246 -422 -244 -397
rect -233 -422 -231 -409
rect -223 -425 -221 -400
rect -216 -425 -214 -400
rect -198 -425 -196 -397
rect -188 -425 -186 -397
rect -178 -425 -176 -397
rect -144 -425 -142 -397
rect -134 -425 -132 -397
rect -124 -425 -122 -397
rect -106 -425 -104 -400
rect -99 -425 -97 -400
rect -89 -422 -87 -409
rect -76 -422 -74 -397
rect 26 -503 28 -475
rect 36 -503 38 -475
rect 46 -503 48 -475
rect 64 -503 66 -478
rect 71 -503 73 -478
rect 81 -500 83 -487
rect 94 -500 96 -475
rect 114 -493 116 -475
rect 121 -493 123 -475
rect 134 -496 136 -484
rect 155 -503 157 -475
rect 165 -503 167 -475
rect 175 -503 177 -475
rect 193 -503 195 -478
rect 200 -503 202 -478
rect 210 -500 212 -487
rect 223 -500 225 -475
rect 245 -500 247 -475
rect 258 -500 260 -487
rect 268 -503 270 -478
rect 275 -503 277 -478
rect 293 -503 295 -475
rect 303 -503 305 -475
rect 313 -503 315 -475
rect 334 -496 336 -484
rect 347 -493 349 -475
rect 354 -493 356 -475
rect 374 -500 376 -475
rect 387 -500 389 -487
rect 397 -503 399 -478
rect 404 -503 406 -478
rect 422 -503 424 -475
rect 432 -503 434 -475
rect 442 -503 444 -475
rect 464 -503 466 -475
rect 474 -503 476 -475
rect 484 -503 486 -475
rect 502 -503 504 -478
rect 509 -503 511 -478
rect 519 -500 521 -487
rect 532 -500 534 -475
rect 552 -493 554 -475
rect 559 -493 561 -475
rect 572 -496 574 -484
rect 593 -503 595 -475
rect 603 -503 605 -475
rect 613 -503 615 -475
rect 631 -503 633 -478
rect 638 -503 640 -478
rect 648 -500 650 -487
rect 661 -500 663 -475
rect 685 -503 687 -475
rect 695 -503 697 -475
rect 705 -503 707 -475
rect 723 -503 725 -478
rect 730 -503 732 -478
rect 740 -500 742 -487
rect 753 -500 755 -475
rect -241 -637 -239 -609
rect -231 -637 -229 -609
rect -221 -637 -219 -609
rect -203 -637 -201 -612
rect -196 -637 -194 -612
rect -186 -634 -184 -621
rect -173 -634 -171 -609
rect -153 -627 -151 -609
rect -146 -627 -144 -609
rect -133 -630 -131 -618
rect -112 -637 -110 -609
rect -102 -637 -100 -609
rect -92 -637 -90 -609
rect -74 -637 -72 -612
rect -67 -637 -65 -612
rect -57 -634 -55 -621
rect -44 -634 -42 -609
rect -22 -634 -20 -609
rect -9 -634 -7 -621
rect 1 -637 3 -612
rect 8 -637 10 -612
rect 26 -637 28 -609
rect 36 -637 38 -609
rect 46 -637 48 -609
rect 67 -630 69 -618
rect 80 -627 82 -609
rect 87 -627 89 -609
rect 107 -634 109 -609
rect 120 -634 122 -621
rect 130 -637 132 -612
rect 137 -637 139 -612
rect 155 -637 157 -609
rect 165 -637 167 -609
rect 175 -637 177 -609
rect 197 -637 199 -609
rect 207 -637 209 -609
rect 217 -637 219 -609
rect 235 -637 237 -612
rect 242 -637 244 -612
rect 252 -634 254 -621
rect 265 -634 267 -609
rect 285 -627 287 -609
rect 292 -627 294 -609
rect 305 -630 307 -618
rect 326 -637 328 -609
rect 336 -637 338 -609
rect 346 -637 348 -609
rect 364 -637 366 -612
rect 371 -637 373 -612
rect 381 -634 383 -621
rect 394 -634 396 -609
rect 418 -637 420 -609
rect 428 -637 430 -609
rect 438 -637 440 -609
rect 456 -637 458 -612
rect 463 -637 465 -612
rect 473 -634 475 -621
rect 486 -634 488 -609
<< polyct0 >>
rect -244 -84 -242 -82
rect -201 -84 -199 -82
rect -158 -84 -156 -82
rect -115 -84 -113 -82
rect -239 -177 -237 -175
rect -245 -187 -243 -185
rect -189 -180 -187 -178
rect -179 -180 -177 -178
rect -145 -180 -143 -178
rect -135 -180 -133 -178
rect -85 -177 -83 -175
rect -79 -187 -77 -185
rect -243 -336 -241 -334
rect -200 -336 -198 -334
rect -157 -336 -155 -334
rect -114 -336 -112 -334
rect 276 158 278 160
rect 319 158 321 160
rect 362 158 364 160
rect 405 158 407 160
rect 281 65 283 67
rect 275 55 277 57
rect 331 62 333 64
rect 341 62 343 64
rect 375 62 377 64
rect 385 62 387 64
rect 435 65 437 67
rect 441 55 443 57
rect 24 -125 26 -123
rect 34 -125 36 -123
rect 84 -122 86 -120
rect 90 -132 92 -130
rect 130 -124 132 -122
rect 153 -125 155 -123
rect 163 -125 165 -123
rect 213 -122 215 -120
rect 219 -132 221 -130
rect 251 -122 253 -120
rect 245 -132 247 -130
rect 301 -125 303 -123
rect 311 -125 313 -123
rect 334 -124 336 -122
rect 380 -122 382 -120
rect 374 -132 376 -130
rect 430 -125 432 -123
rect 440 -125 442 -123
rect 462 -125 464 -123
rect 472 -125 474 -123
rect 522 -122 524 -120
rect 528 -132 530 -130
rect 568 -124 570 -122
rect 591 -125 593 -123
rect 601 -125 603 -123
rect 651 -122 653 -120
rect 683 -125 685 -123
rect 693 -125 695 -123
rect 657 -132 659 -130
rect 743 -122 745 -120
rect 749 -132 751 -130
rect 409 -259 411 -257
rect 452 -259 454 -257
rect 495 -259 497 -257
rect 538 -259 540 -257
rect 414 -352 416 -350
rect 408 -362 410 -360
rect 464 -355 466 -353
rect 474 -355 476 -353
rect 508 -355 510 -353
rect 518 -355 520 -353
rect 568 -352 570 -350
rect 574 -362 576 -360
rect -238 -429 -236 -427
rect -244 -439 -242 -437
rect -188 -432 -186 -430
rect -178 -432 -176 -430
rect -144 -432 -142 -430
rect -134 -432 -132 -430
rect -84 -429 -82 -427
rect -78 -439 -76 -437
rect 26 -510 28 -508
rect 36 -510 38 -508
rect 86 -507 88 -505
rect 92 -517 94 -515
rect 132 -509 134 -507
rect 155 -510 157 -508
rect 165 -510 167 -508
rect 215 -507 217 -505
rect 221 -517 223 -515
rect 253 -507 255 -505
rect 247 -517 249 -515
rect 303 -510 305 -508
rect 313 -510 315 -508
rect 336 -509 338 -507
rect 382 -507 384 -505
rect 376 -517 378 -515
rect 432 -510 434 -508
rect 442 -510 444 -508
rect 464 -510 466 -508
rect 474 -510 476 -508
rect 524 -507 526 -505
rect 530 -517 532 -515
rect 570 -509 572 -507
rect 593 -510 595 -508
rect 603 -510 605 -508
rect 653 -507 655 -505
rect 685 -510 687 -508
rect 695 -510 697 -508
rect 659 -517 661 -515
rect 745 -507 747 -505
rect 751 -517 753 -515
rect -241 -644 -239 -642
rect -231 -644 -229 -642
rect -181 -641 -179 -639
rect -175 -651 -173 -649
rect -135 -643 -133 -641
rect -112 -644 -110 -642
rect -102 -644 -100 -642
rect -52 -641 -50 -639
rect -46 -651 -44 -649
rect -14 -641 -12 -639
rect -20 -651 -18 -649
rect 36 -644 38 -642
rect 46 -644 48 -642
rect 69 -643 71 -641
rect 115 -641 117 -639
rect 109 -651 111 -649
rect 165 -644 167 -642
rect 175 -644 177 -642
rect 197 -644 199 -642
rect 207 -644 209 -642
rect 257 -641 259 -639
rect 263 -651 265 -649
rect 303 -643 305 -641
rect 326 -644 328 -642
rect 336 -644 338 -642
rect 386 -641 388 -639
rect 418 -644 420 -642
rect 428 -644 430 -642
rect 392 -651 394 -649
rect 478 -641 480 -639
rect 484 -651 486 -649
<< polyct1 >>
rect -234 -60 -232 -58
rect -191 -60 -189 -58
rect -105 -60 -103 -58
rect -225 -92 -223 -90
rect -182 -92 -180 -90
rect -139 -92 -137 -90
rect -96 -92 -94 -90
rect -225 -180 -223 -178
rect -206 -180 -204 -178
rect -199 -180 -197 -178
rect -125 -180 -123 -178
rect -118 -180 -116 -178
rect -99 -180 -97 -178
rect -233 -312 -231 -310
rect -190 -312 -188 -310
rect -104 -312 -102 -310
rect -224 -344 -222 -342
rect -181 -344 -179 -342
rect -138 -344 -136 -342
rect -95 -344 -93 -342
rect 286 182 288 184
rect 329 182 331 184
rect 415 182 417 184
rect 295 150 297 152
rect 338 150 340 152
rect 381 150 383 152
rect 424 150 426 152
rect 295 62 297 64
rect 314 62 316 64
rect 321 62 323 64
rect 395 62 397 64
rect 402 62 404 64
rect 421 62 423 64
rect 44 -125 46 -123
rect 51 -125 53 -123
rect 70 -125 72 -123
rect 120 -117 122 -115
rect 110 -125 112 -123
rect 173 -125 175 -123
rect 180 -125 182 -123
rect 199 -125 201 -123
rect 344 -117 346 -115
rect 265 -125 267 -123
rect 284 -125 286 -123
rect 291 -125 293 -123
rect 354 -125 356 -123
rect 394 -125 396 -123
rect 413 -125 415 -123
rect 420 -125 422 -123
rect 482 -125 484 -123
rect 489 -125 491 -123
rect 508 -125 510 -123
rect 558 -117 560 -115
rect 548 -125 550 -123
rect 611 -125 613 -123
rect 618 -125 620 -123
rect 637 -125 639 -123
rect 703 -125 705 -123
rect 710 -125 712 -123
rect 729 -125 731 -123
rect 419 -235 421 -233
rect 462 -235 464 -233
rect 548 -235 550 -233
rect 428 -267 430 -265
rect 471 -267 473 -265
rect 514 -267 516 -265
rect 557 -267 559 -265
rect 591 -308 593 -306
rect 428 -355 430 -353
rect 447 -355 449 -353
rect 454 -355 456 -353
rect 528 -355 530 -353
rect 535 -355 537 -353
rect 554 -355 556 -353
rect -224 -432 -222 -430
rect -205 -432 -203 -430
rect -198 -432 -196 -430
rect -124 -432 -122 -430
rect -117 -432 -115 -430
rect -98 -432 -96 -430
rect 46 -510 48 -508
rect 53 -510 55 -508
rect 72 -510 74 -508
rect 122 -502 124 -500
rect 112 -510 114 -508
rect 175 -510 177 -508
rect 182 -510 184 -508
rect 201 -510 203 -508
rect 346 -502 348 -500
rect 267 -510 269 -508
rect 286 -510 288 -508
rect 293 -510 295 -508
rect 356 -510 358 -508
rect 396 -510 398 -508
rect 415 -510 417 -508
rect 422 -510 424 -508
rect 484 -510 486 -508
rect 491 -510 493 -508
rect 510 -510 512 -508
rect 560 -502 562 -500
rect 550 -510 552 -508
rect 613 -510 615 -508
rect 620 -510 622 -508
rect 639 -510 641 -508
rect 705 -510 707 -508
rect 712 -510 714 -508
rect 731 -510 733 -508
rect -221 -644 -219 -642
rect -214 -644 -212 -642
rect -195 -644 -193 -642
rect -145 -636 -143 -634
rect -155 -644 -153 -642
rect -92 -644 -90 -642
rect -85 -644 -83 -642
rect -66 -644 -64 -642
rect 79 -636 81 -634
rect 0 -644 2 -642
rect 19 -644 21 -642
rect 26 -644 28 -642
rect 89 -644 91 -642
rect 129 -644 131 -642
rect 148 -644 150 -642
rect 155 -644 157 -642
rect 217 -644 219 -642
rect 224 -644 226 -642
rect 243 -644 245 -642
rect 293 -636 295 -634
rect 283 -644 285 -642
rect 346 -644 348 -642
rect 353 -644 355 -642
rect 372 -644 374 -642
rect 438 -644 440 -642
rect 445 -644 447 -642
rect 464 -644 466 -642
<< ndifct0 >>
rect -222 -101 -220 -99
rect -179 -101 -177 -99
rect -136 -101 -134 -99
rect -93 -101 -91 -99
rect -242 -200 -240 -198
rect -232 -197 -230 -195
rect -222 -189 -220 -187
rect -212 -189 -210 -187
rect -212 -196 -210 -194
rect -202 -196 -200 -194
rect -185 -203 -183 -201
rect -139 -203 -137 -201
rect -112 -189 -110 -187
rect -122 -196 -120 -194
rect -112 -196 -110 -194
rect -102 -189 -100 -187
rect -92 -197 -90 -195
rect -82 -200 -80 -198
rect -221 -353 -219 -351
rect -178 -353 -176 -351
rect -135 -353 -133 -351
rect -92 -353 -90 -351
rect 298 141 300 143
rect 341 141 343 143
rect 384 141 386 143
rect 427 141 429 143
rect 278 42 280 44
rect 288 45 290 47
rect 298 53 300 55
rect 308 53 310 55
rect 308 46 310 48
rect 318 46 320 48
rect 335 39 337 41
rect 381 39 383 41
rect 408 53 410 55
rect 398 46 400 48
rect 408 46 410 48
rect 418 53 420 55
rect 428 45 430 47
rect 438 42 440 44
rect 30 -148 32 -146
rect 57 -134 59 -132
rect 47 -141 49 -139
rect 57 -141 59 -139
rect 67 -134 69 -132
rect 77 -142 79 -140
rect 87 -145 89 -143
rect 107 -139 109 -137
rect 117 -139 119 -137
rect 127 -139 129 -137
rect 159 -148 161 -146
rect 186 -134 188 -132
rect 176 -141 178 -139
rect 186 -141 188 -139
rect 196 -134 198 -132
rect 206 -142 208 -140
rect 216 -145 218 -143
rect 248 -145 250 -143
rect 258 -142 260 -140
rect 268 -134 270 -132
rect 278 -134 280 -132
rect 278 -141 280 -139
rect 288 -141 290 -139
rect 305 -148 307 -146
rect 337 -139 339 -137
rect 347 -139 349 -137
rect 357 -139 359 -137
rect 377 -145 379 -143
rect 387 -142 389 -140
rect 397 -134 399 -132
rect 407 -134 409 -132
rect 407 -141 409 -139
rect 417 -141 419 -139
rect 434 -148 436 -146
rect 468 -148 470 -146
rect 495 -134 497 -132
rect 485 -141 487 -139
rect 495 -141 497 -139
rect 505 -134 507 -132
rect 515 -142 517 -140
rect 525 -145 527 -143
rect 545 -139 547 -137
rect 555 -139 557 -137
rect 565 -139 567 -137
rect 597 -148 599 -146
rect 624 -134 626 -132
rect 614 -141 616 -139
rect 624 -141 626 -139
rect 634 -134 636 -132
rect 644 -142 646 -140
rect 654 -145 656 -143
rect 689 -148 691 -146
rect 716 -134 718 -132
rect 706 -141 708 -139
rect 716 -141 718 -139
rect 726 -134 728 -132
rect 736 -142 738 -140
rect 746 -145 748 -143
rect 431 -276 433 -274
rect 474 -276 476 -274
rect 517 -276 519 -274
rect 560 -276 562 -274
rect 411 -375 413 -373
rect 421 -372 423 -370
rect 431 -364 433 -362
rect 441 -364 443 -362
rect 441 -371 443 -369
rect 451 -371 453 -369
rect 468 -378 470 -376
rect 514 -378 516 -376
rect 541 -364 543 -362
rect 531 -371 533 -369
rect 541 -371 543 -369
rect 551 -364 553 -362
rect 561 -372 563 -370
rect 571 -375 573 -373
rect -241 -452 -239 -450
rect -231 -449 -229 -447
rect -221 -441 -219 -439
rect -211 -441 -209 -439
rect -211 -448 -209 -446
rect -201 -448 -199 -446
rect -184 -455 -182 -453
rect -138 -455 -136 -453
rect -111 -441 -109 -439
rect -121 -448 -119 -446
rect -111 -448 -109 -446
rect -101 -441 -99 -439
rect -91 -449 -89 -447
rect -81 -452 -79 -450
rect 32 -533 34 -531
rect 59 -519 61 -517
rect 49 -526 51 -524
rect 59 -526 61 -524
rect 69 -519 71 -517
rect 79 -527 81 -525
rect 89 -530 91 -528
rect 109 -524 111 -522
rect 119 -524 121 -522
rect 129 -524 131 -522
rect 161 -533 163 -531
rect 188 -519 190 -517
rect 178 -526 180 -524
rect 188 -526 190 -524
rect 198 -519 200 -517
rect 208 -527 210 -525
rect 218 -530 220 -528
rect 250 -530 252 -528
rect 260 -527 262 -525
rect 270 -519 272 -517
rect 280 -519 282 -517
rect 280 -526 282 -524
rect 290 -526 292 -524
rect 307 -533 309 -531
rect 339 -524 341 -522
rect 349 -524 351 -522
rect 359 -524 361 -522
rect 379 -530 381 -528
rect 389 -527 391 -525
rect 399 -519 401 -517
rect 409 -519 411 -517
rect 409 -526 411 -524
rect 419 -526 421 -524
rect 436 -533 438 -531
rect 470 -533 472 -531
rect 497 -519 499 -517
rect 487 -526 489 -524
rect 497 -526 499 -524
rect 507 -519 509 -517
rect 517 -527 519 -525
rect 527 -530 529 -528
rect 547 -524 549 -522
rect 557 -524 559 -522
rect 567 -524 569 -522
rect 599 -533 601 -531
rect 626 -519 628 -517
rect 616 -526 618 -524
rect 626 -526 628 -524
rect 636 -519 638 -517
rect 646 -527 648 -525
rect 656 -530 658 -528
rect 691 -533 693 -531
rect 718 -519 720 -517
rect 708 -526 710 -524
rect 718 -526 720 -524
rect 728 -519 730 -517
rect 738 -527 740 -525
rect 748 -530 750 -528
rect -235 -667 -233 -665
rect -208 -653 -206 -651
rect -218 -660 -216 -658
rect -208 -660 -206 -658
rect -198 -653 -196 -651
rect -188 -661 -186 -659
rect -178 -664 -176 -662
rect -158 -658 -156 -656
rect -148 -658 -146 -656
rect -138 -658 -136 -656
rect -106 -667 -104 -665
rect -79 -653 -77 -651
rect -89 -660 -87 -658
rect -79 -660 -77 -658
rect -69 -653 -67 -651
rect -59 -661 -57 -659
rect -49 -664 -47 -662
rect -17 -664 -15 -662
rect -7 -661 -5 -659
rect 3 -653 5 -651
rect 13 -653 15 -651
rect 13 -660 15 -658
rect 23 -660 25 -658
rect 40 -667 42 -665
rect 72 -658 74 -656
rect 82 -658 84 -656
rect 92 -658 94 -656
rect 112 -664 114 -662
rect 122 -661 124 -659
rect 132 -653 134 -651
rect 142 -653 144 -651
rect 142 -660 144 -658
rect 152 -660 154 -658
rect 169 -667 171 -665
rect 203 -667 205 -665
rect 230 -653 232 -651
rect 220 -660 222 -658
rect 230 -660 232 -658
rect 240 -653 242 -651
rect 250 -661 252 -659
rect 260 -664 262 -662
rect 280 -658 282 -656
rect 290 -658 292 -656
rect 300 -658 302 -656
rect 332 -667 334 -665
rect 359 -653 361 -651
rect 349 -660 351 -658
rect 359 -660 361 -658
rect 369 -653 371 -651
rect 379 -661 381 -659
rect 389 -664 391 -662
rect 424 -667 426 -665
rect 451 -653 453 -651
rect 441 -660 443 -658
rect 451 -660 453 -658
rect 461 -653 463 -651
rect 471 -661 473 -659
rect 481 -664 483 -662
<< ndifct1 >>
rect -251 -98 -249 -96
rect -208 -98 -206 -96
rect -165 -98 -163 -96
rect -122 -98 -120 -96
rect -240 -110 -238 -108
rect -197 -110 -195 -108
rect -154 -110 -152 -108
rect -111 -110 -109 -108
rect -252 -196 -250 -194
rect -174 -196 -172 -194
rect -150 -196 -148 -194
rect -72 -196 -70 -194
rect -250 -350 -248 -348
rect -207 -350 -205 -348
rect -164 -350 -162 -348
rect -121 -350 -119 -348
rect -239 -362 -237 -360
rect -196 -362 -194 -360
rect -153 -362 -151 -360
rect -110 -362 -108 -360
rect 269 144 271 146
rect 312 144 314 146
rect 355 144 357 146
rect 398 144 400 146
rect 280 132 282 134
rect 323 132 325 134
rect 366 132 368 134
rect 409 132 411 134
rect 268 46 270 48
rect 346 46 348 48
rect 370 46 372 48
rect 448 46 450 48
rect 19 -141 21 -139
rect 97 -141 99 -139
rect 137 -139 139 -137
rect 148 -141 150 -139
rect 226 -141 228 -139
rect 238 -141 240 -139
rect 316 -141 318 -139
rect 327 -139 329 -137
rect 367 -141 369 -139
rect 445 -141 447 -139
rect 457 -141 459 -139
rect 535 -141 537 -139
rect 575 -139 577 -137
rect 586 -141 588 -139
rect 664 -141 666 -139
rect 678 -141 680 -139
rect 756 -141 758 -139
rect 402 -273 404 -271
rect 445 -273 447 -271
rect 488 -273 490 -271
rect 531 -273 533 -271
rect 413 -285 415 -283
rect 456 -285 458 -283
rect 499 -285 501 -283
rect 542 -285 544 -283
rect 401 -371 403 -369
rect 479 -371 481 -369
rect 503 -371 505 -369
rect 581 -371 583 -369
rect -251 -448 -249 -446
rect -173 -448 -171 -446
rect -149 -448 -147 -446
rect -71 -448 -69 -446
rect 21 -526 23 -524
rect 99 -526 101 -524
rect 139 -524 141 -522
rect 150 -526 152 -524
rect 228 -526 230 -524
rect 240 -526 242 -524
rect 318 -526 320 -524
rect 329 -524 331 -522
rect 369 -526 371 -524
rect 447 -526 449 -524
rect 459 -526 461 -524
rect 537 -526 539 -524
rect 577 -524 579 -522
rect 588 -526 590 -524
rect 666 -526 668 -524
rect 680 -526 682 -524
rect 758 -526 760 -524
rect -246 -660 -244 -658
rect -168 -660 -166 -658
rect -128 -658 -126 -656
rect -117 -660 -115 -658
rect -39 -660 -37 -658
rect -27 -660 -25 -658
rect 51 -660 53 -658
rect 62 -658 64 -656
rect 102 -660 104 -658
rect 180 -660 182 -658
rect 192 -660 194 -658
rect 270 -660 272 -658
rect 310 -658 312 -656
rect 321 -660 323 -658
rect 399 -660 401 -658
rect 413 -660 415 -658
rect 491 -660 493 -658
<< ntiect1 >>
rect 270 192 272 194
rect 284 192 286 194
rect 298 192 300 194
rect 313 192 315 194
rect 327 192 329 194
rect 341 192 343 194
rect 356 192 358 194
rect 370 192 372 194
rect 384 192 386 194
rect 399 192 401 194
rect 413 192 415 194
rect 427 192 429 194
rect -250 -50 -248 -48
rect -236 -50 -234 -48
rect -222 -50 -220 -48
rect -207 -50 -205 -48
rect -193 -50 -191 -48
rect -179 -50 -177 -48
rect -164 -50 -162 -48
rect -150 -50 -148 -48
rect -136 -50 -134 -48
rect -121 -50 -119 -48
rect -107 -50 -105 -48
rect -93 -50 -91 -48
rect -249 -302 -247 -300
rect -235 -302 -233 -300
rect -221 -302 -219 -300
rect -206 -302 -204 -300
rect -192 -302 -190 -300
rect -178 -302 -176 -300
rect -163 -302 -161 -300
rect -149 -302 -147 -300
rect -135 -302 -133 -300
rect -120 -302 -118 -300
rect -106 -302 -104 -300
rect -92 -302 -90 -300
rect 136 -91 138 -89
rect 328 -91 330 -89
rect 574 -91 576 -89
rect 403 -225 405 -223
rect 417 -225 419 -223
rect 431 -225 433 -223
rect 446 -225 448 -223
rect 460 -225 462 -223
rect 474 -225 476 -223
rect 489 -225 491 -223
rect 503 -225 505 -223
rect 517 -225 519 -223
rect 532 -225 534 -223
rect 546 -225 548 -223
rect 560 -225 562 -223
rect 138 -476 140 -474
rect 330 -476 332 -474
rect 576 -476 578 -474
rect -129 -610 -127 -608
rect 63 -610 65 -608
rect 309 -610 311 -608
<< ptiect1 >>
rect -250 -110 -248 -108
rect -207 -110 -205 -108
rect -164 -110 -162 -108
rect -121 -110 -119 -108
rect -249 -362 -247 -360
rect -206 -362 -204 -360
rect -163 -362 -161 -360
rect -120 -362 -118 -360
rect 270 132 272 134
rect 313 132 315 134
rect 356 132 358 134
rect 399 132 401 134
rect 108 -151 110 -149
rect 136 -151 138 -149
rect 328 -151 330 -149
rect 356 -151 358 -149
rect 546 -151 548 -149
rect 574 -151 576 -149
rect 403 -285 405 -283
rect 446 -285 448 -283
rect 489 -285 491 -283
rect 532 -285 534 -283
rect 110 -536 112 -534
rect 138 -536 140 -534
rect 330 -536 332 -534
rect 358 -536 360 -534
rect 548 -536 550 -534
rect 576 -536 578 -534
rect -157 -670 -155 -668
rect -129 -670 -127 -668
rect 63 -670 65 -668
rect 91 -670 93 -668
rect 281 -670 283 -668
rect 309 -670 311 -668
<< pdifct0 >>
rect -241 -75 -239 -73
rect -231 -75 -229 -73
rect -221 -71 -219 -69
rect -198 -75 -196 -73
rect -188 -75 -186 -73
rect -178 -71 -176 -69
rect -155 -75 -153 -73
rect -145 -75 -143 -73
rect -135 -71 -133 -69
rect -112 -75 -110 -73
rect -102 -75 -100 -73
rect -92 -71 -90 -69
rect -241 -149 -239 -147
rect -229 -168 -227 -166
rect -206 -149 -204 -147
rect -206 -156 -204 -154
rect -194 -157 -192 -155
rect -194 -164 -192 -162
rect -184 -149 -182 -147
rect -184 -156 -182 -154
rect -140 -149 -138 -147
rect -140 -156 -138 -154
rect -130 -157 -128 -155
rect -130 -164 -128 -162
rect -118 -149 -116 -147
rect -118 -156 -116 -154
rect -83 -149 -81 -147
rect -95 -168 -93 -166
rect -240 -327 -238 -325
rect -230 -327 -228 -325
rect -220 -323 -218 -321
rect -197 -327 -195 -325
rect -187 -327 -185 -325
rect -177 -323 -175 -321
rect -154 -327 -152 -325
rect -144 -327 -142 -325
rect -134 -323 -132 -321
rect -111 -327 -109 -325
rect -101 -327 -99 -325
rect -91 -323 -89 -321
rect 279 167 281 169
rect 289 167 291 169
rect 299 171 301 173
rect 322 167 324 169
rect 332 167 334 169
rect 342 171 344 173
rect 365 167 367 169
rect 375 167 377 169
rect 385 171 387 173
rect 408 167 410 169
rect 418 167 420 169
rect 428 171 430 173
rect 279 93 281 95
rect 291 74 293 76
rect 314 93 316 95
rect 314 86 316 88
rect 326 85 328 87
rect 326 78 328 80
rect 336 93 338 95
rect 336 86 338 88
rect 380 93 382 95
rect 380 86 382 88
rect 390 85 392 87
rect 390 78 392 80
rect 402 93 404 95
rect 402 86 404 88
rect 437 93 439 95
rect 425 74 427 76
rect 29 -94 31 -92
rect 29 -101 31 -99
rect 39 -102 41 -100
rect 39 -109 41 -107
rect 51 -94 53 -92
rect 51 -101 53 -99
rect 86 -94 88 -92
rect 74 -113 76 -111
rect 107 -101 109 -99
rect 125 -94 127 -92
rect 158 -94 160 -92
rect 158 -101 160 -99
rect 168 -102 170 -100
rect 168 -109 170 -107
rect 180 -94 182 -92
rect 180 -101 182 -99
rect 215 -94 217 -92
rect 203 -113 205 -111
rect 249 -94 251 -92
rect 261 -113 263 -111
rect 284 -94 286 -92
rect 284 -101 286 -99
rect 296 -102 298 -100
rect 296 -109 298 -107
rect 306 -94 308 -92
rect 306 -101 308 -99
rect 339 -94 341 -92
rect 357 -101 359 -99
rect 378 -94 380 -92
rect 390 -113 392 -111
rect 413 -94 415 -92
rect 413 -101 415 -99
rect 425 -102 427 -100
rect 425 -109 427 -107
rect 435 -94 437 -92
rect 435 -101 437 -99
rect 467 -94 469 -92
rect 467 -101 469 -99
rect 477 -102 479 -100
rect 477 -109 479 -107
rect 489 -94 491 -92
rect 489 -101 491 -99
rect 524 -94 526 -92
rect 512 -113 514 -111
rect 545 -101 547 -99
rect 563 -94 565 -92
rect 596 -94 598 -92
rect 596 -101 598 -99
rect 606 -102 608 -100
rect 606 -109 608 -107
rect 618 -94 620 -92
rect 618 -101 620 -99
rect 653 -94 655 -92
rect 641 -113 643 -111
rect 688 -94 690 -92
rect 688 -101 690 -99
rect 698 -102 700 -100
rect 698 -109 700 -107
rect 710 -94 712 -92
rect 710 -101 712 -99
rect 745 -94 747 -92
rect 733 -113 735 -111
rect 412 -250 414 -248
rect 422 -250 424 -248
rect 432 -246 434 -244
rect 455 -250 457 -248
rect 465 -250 467 -248
rect 475 -246 477 -244
rect 498 -250 500 -248
rect 508 -250 510 -248
rect 518 -246 520 -244
rect 541 -250 543 -248
rect 551 -250 553 -248
rect 561 -246 563 -244
rect 412 -324 414 -322
rect 424 -343 426 -341
rect 447 -324 449 -322
rect 447 -331 449 -329
rect 459 -332 461 -330
rect 459 -339 461 -337
rect 469 -324 471 -322
rect 469 -331 471 -329
rect 513 -324 515 -322
rect 513 -331 515 -329
rect 523 -332 525 -330
rect 523 -339 525 -337
rect 535 -324 537 -322
rect 535 -331 537 -329
rect 570 -324 572 -322
rect 558 -343 560 -341
rect -240 -401 -238 -399
rect -228 -420 -226 -418
rect -205 -401 -203 -399
rect -205 -408 -203 -406
rect -193 -409 -191 -407
rect -193 -416 -191 -414
rect -183 -401 -181 -399
rect -183 -408 -181 -406
rect -139 -401 -137 -399
rect -139 -408 -137 -406
rect -129 -409 -127 -407
rect -129 -416 -127 -414
rect -117 -401 -115 -399
rect -117 -408 -115 -406
rect -82 -401 -80 -399
rect -94 -420 -92 -418
rect 31 -479 33 -477
rect 31 -486 33 -484
rect 41 -487 43 -485
rect 41 -494 43 -492
rect 53 -479 55 -477
rect 53 -486 55 -484
rect 88 -479 90 -477
rect 76 -498 78 -496
rect 109 -486 111 -484
rect 127 -479 129 -477
rect 160 -479 162 -477
rect 160 -486 162 -484
rect 170 -487 172 -485
rect 170 -494 172 -492
rect 182 -479 184 -477
rect 182 -486 184 -484
rect 217 -479 219 -477
rect 205 -498 207 -496
rect 251 -479 253 -477
rect 263 -498 265 -496
rect 286 -479 288 -477
rect 286 -486 288 -484
rect 298 -487 300 -485
rect 298 -494 300 -492
rect 308 -479 310 -477
rect 308 -486 310 -484
rect 341 -479 343 -477
rect 359 -486 361 -484
rect 380 -479 382 -477
rect 392 -498 394 -496
rect 415 -479 417 -477
rect 415 -486 417 -484
rect 427 -487 429 -485
rect 427 -494 429 -492
rect 437 -479 439 -477
rect 437 -486 439 -484
rect 469 -479 471 -477
rect 469 -486 471 -484
rect 479 -487 481 -485
rect 479 -494 481 -492
rect 491 -479 493 -477
rect 491 -486 493 -484
rect 526 -479 528 -477
rect 514 -498 516 -496
rect 547 -486 549 -484
rect 565 -479 567 -477
rect 598 -479 600 -477
rect 598 -486 600 -484
rect 608 -487 610 -485
rect 608 -494 610 -492
rect 620 -479 622 -477
rect 620 -486 622 -484
rect 655 -479 657 -477
rect 643 -498 645 -496
rect 690 -479 692 -477
rect 690 -486 692 -484
rect 700 -487 702 -485
rect 700 -494 702 -492
rect 712 -479 714 -477
rect 712 -486 714 -484
rect 747 -479 749 -477
rect 735 -498 737 -496
rect -236 -613 -234 -611
rect -236 -620 -234 -618
rect -226 -621 -224 -619
rect -226 -628 -224 -626
rect -214 -613 -212 -611
rect -214 -620 -212 -618
rect -179 -613 -177 -611
rect -191 -632 -189 -630
rect -158 -620 -156 -618
rect -140 -613 -138 -611
rect -107 -613 -105 -611
rect -107 -620 -105 -618
rect -97 -621 -95 -619
rect -97 -628 -95 -626
rect -85 -613 -83 -611
rect -85 -620 -83 -618
rect -50 -613 -48 -611
rect -62 -632 -60 -630
rect -16 -613 -14 -611
rect -4 -632 -2 -630
rect 19 -613 21 -611
rect 19 -620 21 -618
rect 31 -621 33 -619
rect 31 -628 33 -626
rect 41 -613 43 -611
rect 41 -620 43 -618
rect 74 -613 76 -611
rect 92 -620 94 -618
rect 113 -613 115 -611
rect 125 -632 127 -630
rect 148 -613 150 -611
rect 148 -620 150 -618
rect 160 -621 162 -619
rect 160 -628 162 -626
rect 170 -613 172 -611
rect 170 -620 172 -618
rect 202 -613 204 -611
rect 202 -620 204 -618
rect 212 -621 214 -619
rect 212 -628 214 -626
rect 224 -613 226 -611
rect 224 -620 226 -618
rect 259 -613 261 -611
rect 247 -632 249 -630
rect 280 -620 282 -618
rect 298 -613 300 -611
rect 331 -613 333 -611
rect 331 -620 333 -618
rect 341 -621 343 -619
rect 341 -628 343 -626
rect 353 -613 355 -611
rect 353 -620 355 -618
rect 388 -613 390 -611
rect 376 -632 378 -630
rect 423 -613 425 -611
rect 423 -620 425 -618
rect 433 -621 435 -619
rect 433 -628 435 -626
rect 445 -613 447 -611
rect 445 -620 447 -618
rect 480 -613 482 -611
rect 468 -632 470 -630
<< pdifct1 >>
rect -251 -75 -249 -73
rect -208 -75 -206 -73
rect -165 -75 -163 -73
rect -122 -75 -120 -73
rect -252 -161 -250 -159
rect -252 -168 -250 -166
rect -174 -164 -172 -162
rect -174 -171 -172 -169
rect -150 -164 -148 -162
rect -150 -171 -148 -169
rect -72 -161 -70 -159
rect -72 -168 -70 -166
rect -250 -327 -248 -325
rect -207 -327 -205 -325
rect -164 -327 -162 -325
rect -121 -327 -119 -325
rect 269 167 271 169
rect 312 167 314 169
rect 355 167 357 169
rect 398 167 400 169
rect 268 81 270 83
rect 268 74 270 76
rect 346 78 348 80
rect 346 71 348 73
rect 370 78 372 80
rect 370 71 372 73
rect 448 81 450 83
rect 448 74 450 76
rect 19 -109 21 -107
rect 19 -116 21 -114
rect 97 -106 99 -104
rect 97 -113 99 -111
rect 137 -103 139 -101
rect 148 -109 150 -107
rect 148 -116 150 -114
rect 226 -106 228 -104
rect 226 -113 228 -111
rect 238 -106 240 -104
rect 238 -113 240 -111
rect 327 -103 329 -101
rect 316 -109 318 -107
rect 367 -106 369 -104
rect 316 -116 318 -114
rect 367 -113 369 -111
rect 445 -109 447 -107
rect 445 -116 447 -114
rect 457 -109 459 -107
rect 457 -116 459 -114
rect 535 -106 537 -104
rect 535 -113 537 -111
rect 575 -103 577 -101
rect 586 -109 588 -107
rect 586 -116 588 -114
rect 664 -106 666 -104
rect 664 -113 666 -111
rect 678 -109 680 -107
rect 678 -116 680 -114
rect 756 -106 758 -104
rect 756 -113 758 -111
rect 402 -250 404 -248
rect 445 -250 447 -248
rect 488 -250 490 -248
rect 531 -250 533 -248
rect 401 -336 403 -334
rect 401 -343 403 -341
rect 479 -339 481 -337
rect 479 -346 481 -344
rect 503 -339 505 -337
rect 503 -346 505 -344
rect 581 -336 583 -334
rect 581 -343 583 -341
rect -251 -413 -249 -411
rect -251 -420 -249 -418
rect -173 -416 -171 -414
rect -173 -423 -171 -421
rect -149 -416 -147 -414
rect -149 -423 -147 -421
rect -71 -413 -69 -411
rect -71 -420 -69 -418
rect 21 -494 23 -492
rect 21 -501 23 -499
rect 99 -491 101 -489
rect 99 -498 101 -496
rect 139 -488 141 -486
rect 150 -494 152 -492
rect 150 -501 152 -499
rect 228 -491 230 -489
rect 228 -498 230 -496
rect 240 -491 242 -489
rect 240 -498 242 -496
rect 329 -488 331 -486
rect 318 -494 320 -492
rect 369 -491 371 -489
rect 318 -501 320 -499
rect 369 -498 371 -496
rect 447 -494 449 -492
rect 447 -501 449 -499
rect 459 -494 461 -492
rect 459 -501 461 -499
rect 537 -491 539 -489
rect 537 -498 539 -496
rect 577 -488 579 -486
rect 588 -494 590 -492
rect 588 -501 590 -499
rect 666 -491 668 -489
rect 666 -498 668 -496
rect 680 -494 682 -492
rect 680 -501 682 -499
rect 758 -491 760 -489
rect 758 -498 760 -496
rect -246 -628 -244 -626
rect -246 -635 -244 -633
rect -168 -625 -166 -623
rect -168 -632 -166 -630
rect -128 -622 -126 -620
rect -117 -628 -115 -626
rect -117 -635 -115 -633
rect -39 -625 -37 -623
rect -39 -632 -37 -630
rect -27 -625 -25 -623
rect -27 -632 -25 -630
rect 62 -622 64 -620
rect 51 -628 53 -626
rect 102 -625 104 -623
rect 51 -635 53 -633
rect 102 -632 104 -630
rect 180 -628 182 -626
rect 180 -635 182 -633
rect 192 -628 194 -626
rect 192 -635 194 -633
rect 270 -625 272 -623
rect 270 -632 272 -630
rect 310 -622 312 -620
rect 321 -628 323 -626
rect 321 -635 323 -633
rect 399 -625 401 -623
rect 399 -632 401 -630
rect 413 -628 415 -626
rect 413 -635 415 -633
rect 491 -625 493 -623
rect 491 -632 493 -630
<< alu0 >>
rect 271 165 272 171
rect 275 170 279 191
rect 298 173 302 191
rect 298 171 299 173
rect 301 171 302 173
rect 275 169 283 170
rect 275 167 279 169
rect 281 167 283 169
rect 275 166 283 167
rect 287 169 293 170
rect 298 169 302 171
rect 287 167 289 169
rect 291 167 293 169
rect 287 161 293 167
rect 274 160 293 161
rect 274 158 276 160
rect 278 158 293 160
rect 274 157 293 158
rect 271 146 272 148
rect 283 144 287 157
rect 314 165 315 171
rect 318 170 322 191
rect 341 173 345 191
rect 341 171 342 173
rect 344 171 345 173
rect 318 169 326 170
rect 318 167 322 169
rect 324 167 326 169
rect 318 166 326 167
rect 330 169 336 170
rect 341 169 345 171
rect 330 167 332 169
rect 334 167 336 169
rect 330 161 336 167
rect 317 160 336 161
rect 317 158 319 160
rect 321 158 336 160
rect 317 157 336 158
rect 314 146 315 148
rect 283 143 302 144
rect 283 141 298 143
rect 300 141 302 143
rect 283 140 302 141
rect 326 144 330 157
rect 357 165 358 171
rect 361 170 365 191
rect 384 173 388 191
rect 384 171 385 173
rect 387 171 388 173
rect 361 169 369 170
rect 361 167 365 169
rect 367 167 369 169
rect 361 166 369 167
rect 373 169 379 170
rect 384 169 388 171
rect 373 167 375 169
rect 377 167 379 169
rect 373 161 379 167
rect 360 160 379 161
rect 360 158 362 160
rect 364 158 379 160
rect 360 157 379 158
rect 357 146 358 148
rect 326 143 345 144
rect 326 141 341 143
rect 343 141 345 143
rect 326 140 345 141
rect 369 144 373 157
rect 400 165 401 171
rect 404 170 408 191
rect 427 173 431 191
rect 427 171 428 173
rect 430 171 431 173
rect 404 169 412 170
rect 404 167 408 169
rect 410 167 412 169
rect 404 166 412 167
rect 416 169 422 170
rect 427 169 431 171
rect 416 167 418 169
rect 420 167 422 169
rect 416 161 422 167
rect 403 160 422 161
rect 403 158 405 160
rect 407 158 422 160
rect 403 157 422 158
rect 400 146 401 148
rect 369 143 388 144
rect 369 141 384 143
rect 386 141 388 143
rect 369 140 388 141
rect 412 144 416 157
rect 412 143 431 144
rect 412 141 427 143
rect 429 141 431 143
rect 412 140 431 141
rect 277 93 279 95
rect 281 93 283 95
rect 277 92 283 93
rect 312 93 314 95
rect 316 93 318 95
rect 312 88 318 93
rect 334 93 336 95
rect 338 93 340 95
rect 312 86 314 88
rect 316 86 318 88
rect 312 85 318 86
rect 325 87 329 89
rect 325 85 326 87
rect 328 85 329 87
rect 334 88 340 93
rect 334 86 336 88
rect 338 86 340 88
rect 334 85 340 86
rect 378 93 380 95
rect 382 93 384 95
rect 378 88 384 93
rect 400 93 402 95
rect 404 93 406 95
rect 378 86 380 88
rect 382 86 384 88
rect 378 85 384 86
rect 389 87 393 89
rect 389 85 390 87
rect 392 85 393 87
rect 400 88 406 93
rect 435 93 437 95
rect 439 93 441 95
rect 435 92 441 93
rect 400 86 402 88
rect 404 86 406 88
rect 400 85 406 86
rect 282 81 306 85
rect 325 81 329 85
rect 280 77 286 81
rect 302 80 342 81
rect 302 78 326 80
rect 328 78 342 80
rect 280 67 284 77
rect 290 76 294 78
rect 302 77 342 78
rect 290 74 291 76
rect 293 74 294 76
rect 290 73 294 74
rect 280 65 281 67
rect 283 65 284 67
rect 280 63 284 65
rect 287 69 294 73
rect 287 58 291 69
rect 330 64 334 69
rect 330 62 331 64
rect 333 62 334 64
rect 330 60 334 62
rect 338 66 342 77
rect 338 64 344 66
rect 338 62 341 64
rect 343 62 344 64
rect 338 60 344 62
rect 273 57 291 58
rect 273 55 275 57
rect 277 56 291 57
rect 277 55 302 56
rect 273 54 298 55
rect 287 53 298 54
rect 300 53 302 55
rect 287 52 302 53
rect 307 55 311 57
rect 307 53 308 55
rect 310 53 311 55
rect 307 48 311 53
rect 338 57 342 60
rect 322 53 342 57
rect 389 81 393 85
rect 412 81 436 85
rect 376 80 416 81
rect 376 78 390 80
rect 392 78 416 80
rect 376 77 416 78
rect 376 66 380 77
rect 424 76 428 78
rect 432 77 438 81
rect 424 74 425 76
rect 427 74 428 76
rect 424 73 428 74
rect 424 69 431 73
rect 374 64 380 66
rect 374 62 375 64
rect 377 62 380 64
rect 374 60 380 62
rect 384 64 388 69
rect 384 62 385 64
rect 387 62 388 64
rect 384 60 388 62
rect 322 49 326 53
rect 376 57 380 60
rect 376 53 396 57
rect 392 49 396 53
rect 427 58 431 69
rect 434 67 438 77
rect 434 65 435 67
rect 437 65 438 67
rect 434 63 438 65
rect 427 57 445 58
rect 407 55 411 57
rect 427 56 441 57
rect 407 53 408 55
rect 410 53 411 55
rect 286 47 308 48
rect 277 44 281 46
rect 286 45 288 47
rect 290 46 308 47
rect 310 46 311 48
rect 290 45 311 46
rect 316 48 326 49
rect 316 46 318 48
rect 320 46 326 48
rect 316 45 326 46
rect 392 48 402 49
rect 392 46 398 48
rect 400 46 402 48
rect 392 45 402 46
rect 407 48 411 53
rect 416 55 441 56
rect 443 55 445 57
rect 416 53 418 55
rect 420 54 445 55
rect 420 53 431 54
rect 416 52 431 53
rect 407 46 408 48
rect 410 47 432 48
rect 410 46 428 47
rect 407 45 428 46
rect 430 45 432 47
rect 286 44 311 45
rect 407 44 432 45
rect 437 44 441 46
rect 277 42 278 44
rect 280 42 281 44
rect 437 42 438 44
rect 440 42 441 44
rect 277 39 281 42
rect 333 41 339 42
rect 333 39 335 41
rect 337 39 339 41
rect 379 41 385 42
rect 379 39 381 41
rect 383 39 385 41
rect 437 39 441 42
rect -249 -77 -248 -71
rect -245 -72 -241 -51
rect -222 -69 -218 -51
rect -222 -71 -221 -69
rect -219 -71 -218 -69
rect -245 -73 -237 -72
rect -245 -75 -241 -73
rect -239 -75 -237 -73
rect -245 -76 -237 -75
rect -233 -73 -227 -72
rect -222 -73 -218 -71
rect -233 -75 -231 -73
rect -229 -75 -227 -73
rect -233 -81 -227 -75
rect -246 -82 -227 -81
rect -246 -84 -244 -82
rect -242 -84 -227 -82
rect -246 -85 -227 -84
rect -249 -96 -248 -94
rect -237 -98 -233 -85
rect -206 -77 -205 -71
rect -202 -72 -198 -51
rect -179 -69 -175 -51
rect -179 -71 -178 -69
rect -176 -71 -175 -69
rect -202 -73 -194 -72
rect -202 -75 -198 -73
rect -196 -75 -194 -73
rect -202 -76 -194 -75
rect -190 -73 -184 -72
rect -179 -73 -175 -71
rect -190 -75 -188 -73
rect -186 -75 -184 -73
rect -190 -81 -184 -75
rect -203 -82 -184 -81
rect -203 -84 -201 -82
rect -199 -84 -184 -82
rect -203 -85 -184 -84
rect -206 -96 -205 -94
rect -237 -99 -218 -98
rect -237 -101 -222 -99
rect -220 -101 -218 -99
rect -237 -102 -218 -101
rect -194 -98 -190 -85
rect -163 -77 -162 -71
rect -159 -72 -155 -51
rect -136 -69 -132 -51
rect -136 -71 -135 -69
rect -133 -71 -132 -69
rect -159 -73 -151 -72
rect -159 -75 -155 -73
rect -153 -75 -151 -73
rect -159 -76 -151 -75
rect -147 -73 -141 -72
rect -136 -73 -132 -71
rect -147 -75 -145 -73
rect -143 -75 -141 -73
rect -147 -81 -141 -75
rect -160 -82 -141 -81
rect -160 -84 -158 -82
rect -156 -84 -141 -82
rect -160 -85 -141 -84
rect -163 -96 -162 -94
rect -194 -99 -175 -98
rect -194 -101 -179 -99
rect -177 -101 -175 -99
rect -194 -102 -175 -101
rect -151 -98 -147 -85
rect -120 -77 -119 -71
rect -116 -72 -112 -51
rect -93 -69 -89 -51
rect -93 -71 -92 -69
rect -90 -71 -89 -69
rect -116 -73 -108 -72
rect -116 -75 -112 -73
rect -110 -75 -108 -73
rect -116 -76 -108 -75
rect -104 -73 -98 -72
rect -93 -73 -89 -71
rect -104 -75 -102 -73
rect -100 -75 -98 -73
rect -104 -81 -98 -75
rect -117 -82 -98 -81
rect -117 -84 -115 -82
rect -113 -84 -98 -82
rect -117 -85 -98 -84
rect -120 -96 -119 -94
rect -151 -99 -132 -98
rect -151 -101 -136 -99
rect -134 -101 -132 -99
rect -151 -102 -132 -101
rect -108 -98 -104 -85
rect -108 -99 -89 -98
rect -108 -101 -93 -99
rect -91 -101 -89 -99
rect -108 -102 -89 -101
rect 27 -94 29 -92
rect 31 -94 33 -92
rect 27 -99 33 -94
rect 49 -94 51 -92
rect 53 -94 55 -92
rect 27 -101 29 -99
rect 31 -101 33 -99
rect 27 -102 33 -101
rect 38 -100 42 -98
rect 38 -102 39 -100
rect 41 -102 42 -100
rect 49 -99 55 -94
rect 84 -94 86 -92
rect 88 -94 90 -92
rect 84 -95 90 -94
rect 123 -94 125 -92
rect 127 -94 129 -92
rect 123 -95 129 -94
rect 156 -94 158 -92
rect 160 -94 162 -92
rect 49 -101 51 -99
rect 53 -101 55 -99
rect 49 -102 55 -101
rect 105 -99 125 -98
rect 105 -101 107 -99
rect 109 -101 125 -99
rect 105 -102 125 -101
rect 38 -106 42 -102
rect 61 -106 85 -102
rect 25 -107 65 -106
rect 25 -109 39 -107
rect 41 -109 65 -107
rect 25 -110 65 -109
rect 25 -121 29 -110
rect 73 -111 77 -109
rect 81 -110 87 -106
rect 73 -113 74 -111
rect 76 -113 77 -111
rect 73 -114 77 -113
rect 73 -118 80 -114
rect 23 -123 29 -121
rect 23 -125 24 -123
rect 26 -125 29 -123
rect 23 -127 29 -125
rect 33 -123 37 -118
rect 33 -125 34 -123
rect 36 -125 37 -123
rect 33 -127 37 -125
rect 25 -130 29 -127
rect 25 -134 45 -130
rect 41 -138 45 -134
rect 76 -129 80 -118
rect 83 -120 87 -110
rect 83 -122 84 -120
rect 86 -122 87 -120
rect 83 -124 87 -122
rect 76 -130 94 -129
rect 56 -132 60 -130
rect 76 -131 90 -130
rect 56 -134 57 -132
rect 59 -134 60 -132
rect 41 -139 51 -138
rect 41 -141 47 -139
rect 49 -141 51 -139
rect 41 -142 51 -141
rect 56 -139 60 -134
rect 65 -132 90 -131
rect 92 -132 94 -130
rect 65 -134 67 -132
rect 69 -133 94 -132
rect 69 -134 80 -133
rect 65 -135 80 -134
rect 121 -106 125 -102
rect 136 -105 137 -102
rect 156 -99 162 -94
rect 178 -94 180 -92
rect 182 -94 184 -92
rect 156 -101 158 -99
rect 160 -101 162 -99
rect 156 -102 162 -101
rect 167 -100 171 -98
rect 167 -102 168 -100
rect 170 -102 171 -100
rect 178 -99 184 -94
rect 213 -94 215 -92
rect 217 -94 219 -92
rect 213 -95 219 -94
rect 247 -94 249 -92
rect 251 -94 253 -92
rect 247 -95 253 -94
rect 282 -94 284 -92
rect 286 -94 288 -92
rect 178 -101 180 -99
rect 182 -101 184 -99
rect 178 -102 184 -101
rect 121 -110 133 -106
rect 129 -122 133 -110
rect 129 -124 130 -122
rect 132 -124 133 -122
rect 129 -129 133 -124
rect 116 -133 133 -129
rect 56 -141 57 -139
rect 59 -140 81 -139
rect 59 -141 77 -140
rect 56 -142 77 -141
rect 79 -142 81 -140
rect 56 -143 81 -142
rect 86 -143 90 -141
rect 105 -137 111 -136
rect 105 -139 107 -137
rect 109 -139 111 -137
rect 86 -145 87 -143
rect 89 -145 90 -143
rect -243 -149 -241 -147
rect -239 -149 -237 -147
rect -243 -150 -237 -149
rect -208 -149 -206 -147
rect -204 -149 -202 -147
rect -208 -154 -202 -149
rect -186 -149 -184 -147
rect -182 -149 -180 -147
rect -208 -156 -206 -154
rect -204 -156 -202 -154
rect -208 -157 -202 -156
rect -195 -155 -191 -153
rect -195 -157 -194 -155
rect -192 -157 -191 -155
rect -186 -154 -180 -149
rect -186 -156 -184 -154
rect -182 -156 -180 -154
rect -186 -157 -180 -156
rect -142 -149 -140 -147
rect -138 -149 -136 -147
rect -142 -154 -136 -149
rect -120 -149 -118 -147
rect -116 -149 -114 -147
rect -142 -156 -140 -154
rect -138 -156 -136 -154
rect -142 -157 -136 -156
rect -131 -155 -127 -153
rect -131 -157 -130 -155
rect -128 -157 -127 -155
rect -120 -154 -114 -149
rect -85 -149 -83 -147
rect -81 -149 -79 -147
rect -85 -150 -79 -149
rect -120 -156 -118 -154
rect -116 -156 -114 -154
rect -120 -157 -114 -156
rect -238 -161 -214 -157
rect -195 -161 -191 -157
rect -240 -165 -234 -161
rect -218 -162 -178 -161
rect -218 -164 -194 -162
rect -192 -164 -178 -162
rect -240 -175 -236 -165
rect -230 -166 -226 -164
rect -218 -165 -178 -164
rect -230 -168 -229 -166
rect -227 -168 -226 -166
rect -230 -169 -226 -168
rect -240 -177 -239 -175
rect -237 -177 -236 -175
rect -240 -179 -236 -177
rect -233 -173 -226 -169
rect -233 -184 -229 -173
rect -190 -178 -186 -173
rect -190 -180 -189 -178
rect -187 -180 -186 -178
rect -190 -182 -186 -180
rect -182 -176 -178 -165
rect -182 -178 -176 -176
rect -182 -180 -179 -178
rect -177 -180 -176 -178
rect -182 -182 -176 -180
rect -247 -185 -229 -184
rect -247 -187 -245 -185
rect -243 -186 -229 -185
rect -243 -187 -218 -186
rect -247 -188 -222 -187
rect -233 -189 -222 -188
rect -220 -189 -218 -187
rect -233 -190 -218 -189
rect -213 -187 -209 -185
rect -213 -189 -212 -187
rect -210 -189 -209 -187
rect -213 -194 -209 -189
rect -182 -185 -178 -182
rect -198 -189 -178 -185
rect -198 -193 -194 -189
rect -131 -161 -127 -157
rect -108 -161 -84 -157
rect -144 -162 -104 -161
rect -144 -164 -130 -162
rect -128 -164 -104 -162
rect -144 -165 -104 -164
rect -144 -176 -140 -165
rect -96 -166 -92 -164
rect -88 -165 -82 -161
rect -96 -168 -95 -166
rect -93 -168 -92 -166
rect -96 -169 -92 -168
rect -96 -173 -89 -169
rect -146 -178 -140 -176
rect -146 -180 -145 -178
rect -143 -180 -140 -178
rect -146 -182 -140 -180
rect -136 -178 -132 -173
rect -136 -180 -135 -178
rect -133 -180 -132 -178
rect -136 -182 -132 -180
rect -234 -195 -212 -194
rect -243 -198 -239 -196
rect -234 -197 -232 -195
rect -230 -196 -212 -195
rect -210 -196 -209 -194
rect -230 -197 -209 -196
rect -204 -194 -194 -193
rect -204 -196 -202 -194
rect -200 -196 -194 -194
rect -204 -197 -194 -196
rect -144 -185 -140 -182
rect -144 -189 -124 -185
rect -128 -193 -124 -189
rect -93 -184 -89 -173
rect -86 -175 -82 -165
rect -86 -177 -85 -175
rect -83 -177 -82 -175
rect -86 -179 -82 -177
rect -93 -185 -75 -184
rect -113 -187 -109 -185
rect -93 -186 -79 -185
rect -113 -189 -112 -187
rect -110 -189 -109 -187
rect -128 -194 -118 -193
rect -128 -196 -122 -194
rect -120 -196 -118 -194
rect -128 -197 -118 -196
rect -113 -194 -109 -189
rect -104 -187 -79 -186
rect -77 -187 -75 -185
rect -104 -189 -102 -187
rect -100 -188 -75 -187
rect -100 -189 -89 -188
rect -104 -190 -89 -189
rect -113 -196 -112 -194
rect -110 -195 -88 -194
rect -110 -196 -92 -195
rect -113 -197 -92 -196
rect -90 -197 -88 -195
rect -234 -198 -209 -197
rect -113 -198 -88 -197
rect -83 -198 -79 -196
rect -243 -200 -242 -198
rect -240 -200 -239 -198
rect -83 -200 -82 -198
rect -80 -200 -79 -198
rect -243 -203 -239 -200
rect -187 -201 -181 -200
rect -187 -203 -185 -201
rect -183 -203 -181 -201
rect -141 -201 -135 -200
rect -141 -203 -139 -201
rect -137 -203 -135 -201
rect -83 -203 -79 -200
rect 28 -146 34 -145
rect 28 -148 30 -146
rect 32 -148 34 -146
rect 86 -148 90 -145
rect 105 -148 111 -139
rect 116 -137 120 -133
rect 116 -139 117 -137
rect 119 -139 120 -137
rect 116 -141 120 -139
rect 125 -137 131 -136
rect 125 -139 127 -137
rect 129 -139 131 -137
rect 125 -148 131 -139
rect 167 -106 171 -102
rect 190 -106 214 -102
rect 154 -107 194 -106
rect 154 -109 168 -107
rect 170 -109 194 -107
rect 154 -110 194 -109
rect 154 -121 158 -110
rect 202 -111 206 -109
rect 210 -110 216 -106
rect 202 -113 203 -111
rect 205 -113 206 -111
rect 202 -114 206 -113
rect 202 -118 209 -114
rect 152 -123 158 -121
rect 152 -125 153 -123
rect 155 -125 158 -123
rect 152 -127 158 -125
rect 162 -123 166 -118
rect 162 -125 163 -123
rect 165 -125 166 -123
rect 162 -127 166 -125
rect 154 -130 158 -127
rect 154 -134 174 -130
rect 170 -138 174 -134
rect 205 -129 209 -118
rect 212 -120 216 -110
rect 212 -122 213 -120
rect 215 -122 216 -120
rect 212 -124 216 -122
rect 205 -130 223 -129
rect 185 -132 189 -130
rect 205 -131 219 -130
rect 185 -134 186 -132
rect 188 -134 189 -132
rect 170 -139 180 -138
rect 170 -141 176 -139
rect 178 -141 180 -139
rect 170 -142 180 -141
rect 185 -139 189 -134
rect 194 -132 219 -131
rect 221 -132 223 -130
rect 194 -134 196 -132
rect 198 -133 223 -132
rect 198 -134 209 -133
rect 194 -135 209 -134
rect 185 -141 186 -139
rect 188 -140 210 -139
rect 188 -141 206 -140
rect 185 -142 206 -141
rect 208 -142 210 -140
rect 185 -143 210 -142
rect 215 -143 219 -141
rect 282 -99 288 -94
rect 304 -94 306 -92
rect 308 -94 310 -92
rect 282 -101 284 -99
rect 286 -101 288 -99
rect 282 -102 288 -101
rect 295 -100 299 -98
rect 295 -102 296 -100
rect 298 -102 299 -100
rect 304 -99 310 -94
rect 337 -94 339 -92
rect 341 -94 343 -92
rect 337 -95 343 -94
rect 376 -94 378 -92
rect 380 -94 382 -92
rect 376 -95 382 -94
rect 411 -94 413 -92
rect 415 -94 417 -92
rect 304 -101 306 -99
rect 308 -101 310 -99
rect 304 -102 310 -101
rect 252 -106 276 -102
rect 295 -106 299 -102
rect 341 -99 361 -98
rect 341 -101 357 -99
rect 359 -101 361 -99
rect 341 -102 361 -101
rect 411 -99 417 -94
rect 433 -94 435 -92
rect 437 -94 439 -92
rect 411 -101 413 -99
rect 415 -101 417 -99
rect 411 -102 417 -101
rect 424 -100 428 -98
rect 424 -102 425 -100
rect 427 -102 428 -100
rect 433 -99 439 -94
rect 433 -101 435 -99
rect 437 -101 439 -99
rect 433 -102 439 -101
rect 465 -94 467 -92
rect 469 -94 471 -92
rect 465 -99 471 -94
rect 487 -94 489 -92
rect 491 -94 493 -92
rect 465 -101 467 -99
rect 469 -101 471 -99
rect 465 -102 471 -101
rect 476 -100 480 -98
rect 476 -102 477 -100
rect 479 -102 480 -100
rect 487 -99 493 -94
rect 522 -94 524 -92
rect 526 -94 528 -92
rect 522 -95 528 -94
rect 561 -94 563 -92
rect 565 -94 567 -92
rect 561 -95 567 -94
rect 594 -94 596 -92
rect 598 -94 600 -92
rect 487 -101 489 -99
rect 491 -101 493 -99
rect 487 -102 493 -101
rect 543 -99 563 -98
rect 543 -101 545 -99
rect 547 -101 563 -99
rect 543 -102 563 -101
rect 250 -110 256 -106
rect 272 -107 312 -106
rect 272 -109 296 -107
rect 298 -109 312 -107
rect 250 -120 254 -110
rect 260 -111 264 -109
rect 272 -110 312 -109
rect 260 -113 261 -111
rect 263 -113 264 -111
rect 260 -114 264 -113
rect 250 -122 251 -120
rect 253 -122 254 -120
rect 250 -124 254 -122
rect 257 -118 264 -114
rect 257 -129 261 -118
rect 300 -123 304 -118
rect 300 -125 301 -123
rect 303 -125 304 -123
rect 243 -130 261 -129
rect 243 -132 245 -130
rect 247 -131 261 -130
rect 247 -132 272 -131
rect 243 -133 268 -132
rect 257 -134 268 -133
rect 270 -134 272 -132
rect 257 -135 272 -134
rect 277 -132 281 -130
rect 277 -134 278 -132
rect 280 -134 281 -132
rect 277 -139 281 -134
rect 300 -127 304 -125
rect 308 -121 312 -110
rect 308 -123 314 -121
rect 308 -125 311 -123
rect 313 -125 314 -123
rect 308 -127 314 -125
rect 308 -130 312 -127
rect 292 -134 312 -130
rect 292 -138 296 -134
rect 256 -140 278 -139
rect 247 -143 251 -141
rect 256 -142 258 -140
rect 260 -141 278 -140
rect 280 -141 281 -139
rect 260 -142 281 -141
rect 286 -139 296 -138
rect 286 -141 288 -139
rect 290 -141 296 -139
rect 286 -142 296 -141
rect 329 -105 330 -102
rect 341 -106 345 -102
rect 333 -110 345 -106
rect 333 -122 337 -110
rect 381 -106 405 -102
rect 424 -106 428 -102
rect 333 -124 334 -122
rect 336 -124 337 -122
rect 333 -129 337 -124
rect 379 -110 385 -106
rect 401 -107 441 -106
rect 401 -109 425 -107
rect 427 -109 441 -107
rect 379 -120 383 -110
rect 389 -111 393 -109
rect 401 -110 441 -109
rect 389 -113 390 -111
rect 392 -113 393 -111
rect 389 -114 393 -113
rect 379 -122 380 -120
rect 382 -122 383 -120
rect 379 -124 383 -122
rect 386 -118 393 -114
rect 333 -133 350 -129
rect 256 -143 281 -142
rect 335 -137 341 -136
rect 335 -139 337 -137
rect 339 -139 341 -137
rect 215 -145 216 -143
rect 218 -145 219 -143
rect 157 -146 163 -145
rect 157 -148 159 -146
rect 161 -148 163 -146
rect 215 -148 219 -145
rect 247 -145 248 -143
rect 250 -145 251 -143
rect 247 -148 251 -145
rect 303 -146 309 -145
rect 303 -148 305 -146
rect 307 -148 309 -146
rect 335 -148 341 -139
rect 346 -137 350 -133
rect 346 -139 347 -137
rect 349 -139 350 -137
rect 346 -141 350 -139
rect 355 -137 361 -136
rect 355 -139 357 -137
rect 359 -139 361 -137
rect 355 -148 361 -139
rect 386 -129 390 -118
rect 429 -123 433 -118
rect 429 -125 430 -123
rect 432 -125 433 -123
rect 372 -130 390 -129
rect 429 -127 433 -125
rect 437 -121 441 -110
rect 437 -123 443 -121
rect 437 -125 440 -123
rect 442 -125 443 -123
rect 437 -127 443 -125
rect 372 -132 374 -130
rect 376 -131 390 -130
rect 376 -132 401 -131
rect 372 -133 397 -132
rect 386 -134 397 -133
rect 399 -134 401 -132
rect 386 -135 401 -134
rect 406 -132 410 -130
rect 406 -134 407 -132
rect 409 -134 410 -132
rect 406 -139 410 -134
rect 437 -130 441 -127
rect 421 -134 441 -130
rect 421 -138 425 -134
rect 385 -140 407 -139
rect 376 -143 380 -141
rect 385 -142 387 -140
rect 389 -141 407 -140
rect 409 -141 410 -139
rect 389 -142 410 -141
rect 415 -139 425 -138
rect 415 -141 417 -139
rect 419 -141 425 -139
rect 415 -142 425 -141
rect 476 -106 480 -102
rect 499 -106 523 -102
rect 463 -107 503 -106
rect 463 -109 477 -107
rect 479 -109 503 -107
rect 463 -110 503 -109
rect 463 -121 467 -110
rect 511 -111 515 -109
rect 519 -110 525 -106
rect 511 -113 512 -111
rect 514 -113 515 -111
rect 511 -114 515 -113
rect 511 -118 518 -114
rect 461 -123 467 -121
rect 461 -125 462 -123
rect 464 -125 467 -123
rect 461 -127 467 -125
rect 471 -123 475 -118
rect 471 -125 472 -123
rect 474 -125 475 -123
rect 471 -127 475 -125
rect 463 -130 467 -127
rect 463 -134 483 -130
rect 479 -138 483 -134
rect 514 -129 518 -118
rect 521 -120 525 -110
rect 521 -122 522 -120
rect 524 -122 525 -120
rect 521 -124 525 -122
rect 514 -130 532 -129
rect 494 -132 498 -130
rect 514 -131 528 -130
rect 494 -134 495 -132
rect 497 -134 498 -132
rect 479 -139 489 -138
rect 479 -141 485 -139
rect 487 -141 489 -139
rect 479 -142 489 -141
rect 494 -139 498 -134
rect 503 -132 528 -131
rect 530 -132 532 -130
rect 503 -134 505 -132
rect 507 -133 532 -132
rect 507 -134 518 -133
rect 503 -135 518 -134
rect 559 -106 563 -102
rect 574 -105 575 -102
rect 594 -99 600 -94
rect 616 -94 618 -92
rect 620 -94 622 -92
rect 594 -101 596 -99
rect 598 -101 600 -99
rect 594 -102 600 -101
rect 605 -100 609 -98
rect 605 -102 606 -100
rect 608 -102 609 -100
rect 616 -99 622 -94
rect 651 -94 653 -92
rect 655 -94 657 -92
rect 651 -95 657 -94
rect 686 -94 688 -92
rect 690 -94 692 -92
rect 616 -101 618 -99
rect 620 -101 622 -99
rect 616 -102 622 -101
rect 686 -99 692 -94
rect 708 -94 710 -92
rect 712 -94 714 -92
rect 686 -101 688 -99
rect 690 -101 692 -99
rect 686 -102 692 -101
rect 697 -100 701 -98
rect 697 -102 698 -100
rect 700 -102 701 -100
rect 708 -99 714 -94
rect 743 -94 745 -92
rect 747 -94 749 -92
rect 743 -95 749 -94
rect 708 -101 710 -99
rect 712 -101 714 -99
rect 708 -102 714 -101
rect 559 -110 571 -106
rect 567 -122 571 -110
rect 567 -124 568 -122
rect 570 -124 571 -122
rect 567 -129 571 -124
rect 554 -133 571 -129
rect 494 -141 495 -139
rect 497 -140 519 -139
rect 497 -141 515 -140
rect 494 -142 515 -141
rect 517 -142 519 -140
rect 385 -143 410 -142
rect 494 -143 519 -142
rect 524 -143 528 -141
rect 543 -137 549 -136
rect 543 -139 545 -137
rect 547 -139 549 -137
rect 376 -145 377 -143
rect 379 -145 380 -143
rect 524 -145 525 -143
rect 527 -145 528 -143
rect 376 -148 380 -145
rect 432 -146 438 -145
rect 432 -148 434 -146
rect 436 -148 438 -146
rect 466 -146 472 -145
rect 466 -148 468 -146
rect 470 -148 472 -146
rect 524 -148 528 -145
rect 543 -148 549 -139
rect 554 -137 558 -133
rect 554 -139 555 -137
rect 557 -139 558 -137
rect 554 -141 558 -139
rect 563 -137 569 -136
rect 563 -139 565 -137
rect 567 -139 569 -137
rect 563 -148 569 -139
rect 605 -106 609 -102
rect 628 -106 652 -102
rect 592 -107 632 -106
rect 592 -109 606 -107
rect 608 -109 632 -107
rect 592 -110 632 -109
rect 592 -121 596 -110
rect 640 -111 644 -109
rect 648 -110 654 -106
rect 640 -113 641 -111
rect 643 -113 644 -111
rect 640 -114 644 -113
rect 640 -118 647 -114
rect 590 -123 596 -121
rect 590 -125 591 -123
rect 593 -125 596 -123
rect 590 -127 596 -125
rect 600 -123 604 -118
rect 600 -125 601 -123
rect 603 -125 604 -123
rect 600 -127 604 -125
rect 592 -130 596 -127
rect 592 -134 612 -130
rect 608 -138 612 -134
rect 643 -129 647 -118
rect 650 -120 654 -110
rect 650 -122 651 -120
rect 653 -122 654 -120
rect 650 -124 654 -122
rect 643 -130 661 -129
rect 623 -132 627 -130
rect 643 -131 657 -130
rect 623 -134 624 -132
rect 626 -134 627 -132
rect 608 -139 618 -138
rect 608 -141 614 -139
rect 616 -141 618 -139
rect 608 -142 618 -141
rect 623 -139 627 -134
rect 632 -132 657 -131
rect 659 -132 661 -130
rect 632 -134 634 -132
rect 636 -133 661 -132
rect 636 -134 647 -133
rect 632 -135 647 -134
rect 623 -141 624 -139
rect 626 -140 648 -139
rect 626 -141 644 -140
rect 623 -142 644 -141
rect 646 -142 648 -140
rect 623 -143 648 -142
rect 653 -143 657 -141
rect 697 -106 701 -102
rect 720 -106 744 -102
rect 684 -107 724 -106
rect 684 -109 698 -107
rect 700 -109 724 -107
rect 684 -110 724 -109
rect 684 -121 688 -110
rect 732 -111 736 -109
rect 740 -110 746 -106
rect 732 -113 733 -111
rect 735 -113 736 -111
rect 732 -114 736 -113
rect 732 -118 739 -114
rect 682 -123 688 -121
rect 682 -125 683 -123
rect 685 -125 688 -123
rect 682 -127 688 -125
rect 692 -123 696 -118
rect 692 -125 693 -123
rect 695 -125 696 -123
rect 692 -127 696 -125
rect 684 -130 688 -127
rect 684 -134 704 -130
rect 700 -138 704 -134
rect 735 -129 739 -118
rect 742 -120 746 -110
rect 742 -122 743 -120
rect 745 -122 746 -120
rect 742 -124 746 -122
rect 735 -130 753 -129
rect 715 -132 719 -130
rect 735 -131 749 -130
rect 715 -134 716 -132
rect 718 -134 719 -132
rect 700 -139 710 -138
rect 700 -141 706 -139
rect 708 -141 710 -139
rect 700 -142 710 -141
rect 715 -139 719 -134
rect 724 -132 749 -131
rect 751 -132 753 -130
rect 724 -134 726 -132
rect 728 -133 753 -132
rect 728 -134 739 -133
rect 724 -135 739 -134
rect 715 -141 716 -139
rect 718 -140 740 -139
rect 718 -141 736 -140
rect 715 -142 736 -141
rect 738 -142 740 -140
rect 715 -143 740 -142
rect 745 -143 749 -141
rect 653 -145 654 -143
rect 656 -145 657 -143
rect 745 -145 746 -143
rect 748 -145 749 -143
rect 595 -146 601 -145
rect 595 -148 597 -146
rect 599 -148 601 -146
rect 653 -148 657 -145
rect 687 -146 693 -145
rect 687 -148 689 -146
rect 691 -148 693 -146
rect 745 -148 749 -145
rect -248 -329 -247 -323
rect -244 -324 -240 -303
rect -221 -321 -217 -303
rect -221 -323 -220 -321
rect -218 -323 -217 -321
rect -244 -325 -236 -324
rect -244 -327 -240 -325
rect -238 -327 -236 -325
rect -244 -328 -236 -327
rect -232 -325 -226 -324
rect -221 -325 -217 -323
rect -232 -327 -230 -325
rect -228 -327 -226 -325
rect -232 -333 -226 -327
rect -245 -334 -226 -333
rect -245 -336 -243 -334
rect -241 -336 -226 -334
rect -245 -337 -226 -336
rect -248 -348 -247 -346
rect -236 -350 -232 -337
rect -205 -329 -204 -323
rect -201 -324 -197 -303
rect -178 -321 -174 -303
rect -178 -323 -177 -321
rect -175 -323 -174 -321
rect -201 -325 -193 -324
rect -201 -327 -197 -325
rect -195 -327 -193 -325
rect -201 -328 -193 -327
rect -189 -325 -183 -324
rect -178 -325 -174 -323
rect -189 -327 -187 -325
rect -185 -327 -183 -325
rect -189 -333 -183 -327
rect -202 -334 -183 -333
rect -202 -336 -200 -334
rect -198 -336 -183 -334
rect -202 -337 -183 -336
rect -205 -348 -204 -346
rect -236 -351 -217 -350
rect -236 -353 -221 -351
rect -219 -353 -217 -351
rect -236 -354 -217 -353
rect -193 -350 -189 -337
rect -162 -329 -161 -323
rect -158 -324 -154 -303
rect -135 -321 -131 -303
rect -135 -323 -134 -321
rect -132 -323 -131 -321
rect -158 -325 -150 -324
rect -158 -327 -154 -325
rect -152 -327 -150 -325
rect -158 -328 -150 -327
rect -146 -325 -140 -324
rect -135 -325 -131 -323
rect -146 -327 -144 -325
rect -142 -327 -140 -325
rect -146 -333 -140 -327
rect -159 -334 -140 -333
rect -159 -336 -157 -334
rect -155 -336 -140 -334
rect -159 -337 -140 -336
rect -162 -348 -161 -346
rect -193 -351 -174 -350
rect -193 -353 -178 -351
rect -176 -353 -174 -351
rect -193 -354 -174 -353
rect -150 -350 -146 -337
rect -119 -329 -118 -323
rect -115 -324 -111 -303
rect -92 -321 -88 -303
rect -92 -323 -91 -321
rect -89 -323 -88 -321
rect -115 -325 -107 -324
rect -115 -327 -111 -325
rect -109 -327 -107 -325
rect -115 -328 -107 -327
rect -103 -325 -97 -324
rect -92 -325 -88 -323
rect -103 -327 -101 -325
rect -99 -327 -97 -325
rect -103 -333 -97 -327
rect -116 -334 -97 -333
rect -116 -336 -114 -334
rect -112 -336 -97 -334
rect -116 -337 -97 -336
rect -119 -348 -118 -346
rect -150 -351 -131 -350
rect -150 -353 -135 -351
rect -133 -353 -131 -351
rect -150 -354 -131 -353
rect -107 -350 -103 -337
rect -107 -351 -88 -350
rect -107 -353 -92 -351
rect -90 -353 -88 -351
rect -107 -354 -88 -353
rect 404 -252 405 -246
rect 408 -247 412 -226
rect 431 -244 435 -226
rect 431 -246 432 -244
rect 434 -246 435 -244
rect 408 -248 416 -247
rect 408 -250 412 -248
rect 414 -250 416 -248
rect 408 -251 416 -250
rect 420 -248 426 -247
rect 431 -248 435 -246
rect 420 -250 422 -248
rect 424 -250 426 -248
rect 420 -256 426 -250
rect 407 -257 426 -256
rect 407 -259 409 -257
rect 411 -259 426 -257
rect 407 -260 426 -259
rect 404 -271 405 -269
rect 416 -273 420 -260
rect 447 -252 448 -246
rect 451 -247 455 -226
rect 474 -244 478 -226
rect 474 -246 475 -244
rect 477 -246 478 -244
rect 451 -248 459 -247
rect 451 -250 455 -248
rect 457 -250 459 -248
rect 451 -251 459 -250
rect 463 -248 469 -247
rect 474 -248 478 -246
rect 463 -250 465 -248
rect 467 -250 469 -248
rect 463 -256 469 -250
rect 450 -257 469 -256
rect 450 -259 452 -257
rect 454 -259 469 -257
rect 450 -260 469 -259
rect 447 -271 448 -269
rect 416 -274 435 -273
rect 416 -276 431 -274
rect 433 -276 435 -274
rect 416 -277 435 -276
rect 459 -273 463 -260
rect 490 -252 491 -246
rect 494 -247 498 -226
rect 517 -244 521 -226
rect 517 -246 518 -244
rect 520 -246 521 -244
rect 494 -248 502 -247
rect 494 -250 498 -248
rect 500 -250 502 -248
rect 494 -251 502 -250
rect 506 -248 512 -247
rect 517 -248 521 -246
rect 506 -250 508 -248
rect 510 -250 512 -248
rect 506 -256 512 -250
rect 493 -257 512 -256
rect 493 -259 495 -257
rect 497 -259 512 -257
rect 493 -260 512 -259
rect 490 -271 491 -269
rect 459 -274 478 -273
rect 459 -276 474 -274
rect 476 -276 478 -274
rect 459 -277 478 -276
rect 502 -273 506 -260
rect 533 -252 534 -246
rect 537 -247 541 -226
rect 560 -244 564 -226
rect 560 -246 561 -244
rect 563 -246 564 -244
rect 537 -248 545 -247
rect 537 -250 541 -248
rect 543 -250 545 -248
rect 537 -251 545 -250
rect 549 -248 555 -247
rect 560 -248 564 -246
rect 549 -250 551 -248
rect 553 -250 555 -248
rect 549 -256 555 -250
rect 536 -257 555 -256
rect 536 -259 538 -257
rect 540 -259 555 -257
rect 536 -260 555 -259
rect 533 -271 534 -269
rect 502 -274 521 -273
rect 502 -276 517 -274
rect 519 -276 521 -274
rect 502 -277 521 -276
rect 545 -273 549 -260
rect 545 -274 564 -273
rect 545 -276 560 -274
rect 562 -276 564 -274
rect 545 -277 564 -276
rect 410 -324 412 -322
rect 414 -324 416 -322
rect 410 -325 416 -324
rect 445 -324 447 -322
rect 449 -324 451 -322
rect 445 -329 451 -324
rect 467 -324 469 -322
rect 471 -324 473 -322
rect 445 -331 447 -329
rect 449 -331 451 -329
rect 445 -332 451 -331
rect 458 -330 462 -328
rect 458 -332 459 -330
rect 461 -332 462 -330
rect 467 -329 473 -324
rect 467 -331 469 -329
rect 471 -331 473 -329
rect 467 -332 473 -331
rect 511 -324 513 -322
rect 515 -324 517 -322
rect 511 -329 517 -324
rect 533 -324 535 -322
rect 537 -324 539 -322
rect 511 -331 513 -329
rect 515 -331 517 -329
rect 511 -332 517 -331
rect 522 -330 526 -328
rect 522 -332 523 -330
rect 525 -332 526 -330
rect 533 -329 539 -324
rect 568 -324 570 -322
rect 572 -324 574 -322
rect 568 -325 574 -324
rect 533 -331 535 -329
rect 537 -331 539 -329
rect 533 -332 539 -331
rect 415 -336 439 -332
rect 458 -336 462 -332
rect 413 -340 419 -336
rect 435 -337 475 -336
rect 435 -339 459 -337
rect 461 -339 475 -337
rect 413 -350 417 -340
rect 423 -341 427 -339
rect 435 -340 475 -339
rect 423 -343 424 -341
rect 426 -343 427 -341
rect 423 -344 427 -343
rect 413 -352 414 -350
rect 416 -352 417 -350
rect 413 -354 417 -352
rect 420 -348 427 -344
rect -242 -401 -240 -399
rect -238 -401 -236 -399
rect -242 -402 -236 -401
rect -207 -401 -205 -399
rect -203 -401 -201 -399
rect -207 -406 -201 -401
rect -185 -401 -183 -399
rect -181 -401 -179 -399
rect -207 -408 -205 -406
rect -203 -408 -201 -406
rect -207 -409 -201 -408
rect -194 -407 -190 -405
rect -194 -409 -193 -407
rect -191 -409 -190 -407
rect -185 -406 -179 -401
rect -185 -408 -183 -406
rect -181 -408 -179 -406
rect -185 -409 -179 -408
rect -141 -401 -139 -399
rect -137 -401 -135 -399
rect -141 -406 -135 -401
rect -119 -401 -117 -399
rect -115 -401 -113 -399
rect -141 -408 -139 -406
rect -137 -408 -135 -406
rect -141 -409 -135 -408
rect -130 -407 -126 -405
rect -130 -409 -129 -407
rect -127 -409 -126 -407
rect -119 -406 -113 -401
rect -84 -401 -82 -399
rect -80 -401 -78 -399
rect -84 -402 -78 -401
rect -119 -408 -117 -406
rect -115 -408 -113 -406
rect -119 -409 -113 -408
rect -237 -413 -213 -409
rect -194 -413 -190 -409
rect -239 -417 -233 -413
rect -217 -414 -177 -413
rect -217 -416 -193 -414
rect -191 -416 -177 -414
rect -239 -427 -235 -417
rect -229 -418 -225 -416
rect -217 -417 -177 -416
rect -229 -420 -228 -418
rect -226 -420 -225 -418
rect -229 -421 -225 -420
rect -239 -429 -238 -427
rect -236 -429 -235 -427
rect -239 -431 -235 -429
rect -232 -425 -225 -421
rect -232 -436 -228 -425
rect -189 -430 -185 -425
rect -189 -432 -188 -430
rect -186 -432 -185 -430
rect -189 -434 -185 -432
rect -181 -428 -177 -417
rect -181 -430 -175 -428
rect -181 -432 -178 -430
rect -176 -432 -175 -430
rect -181 -434 -175 -432
rect -246 -437 -228 -436
rect -246 -439 -244 -437
rect -242 -438 -228 -437
rect -242 -439 -217 -438
rect -246 -440 -221 -439
rect -232 -441 -221 -440
rect -219 -441 -217 -439
rect -232 -442 -217 -441
rect -212 -439 -208 -437
rect -212 -441 -211 -439
rect -209 -441 -208 -439
rect -212 -446 -208 -441
rect -181 -437 -177 -434
rect -197 -441 -177 -437
rect -197 -445 -193 -441
rect -130 -413 -126 -409
rect -107 -413 -83 -409
rect -143 -414 -103 -413
rect -143 -416 -129 -414
rect -127 -416 -103 -414
rect -143 -417 -103 -416
rect -143 -428 -139 -417
rect -95 -418 -91 -416
rect -87 -417 -81 -413
rect -95 -420 -94 -418
rect -92 -420 -91 -418
rect -95 -421 -91 -420
rect -95 -425 -88 -421
rect -145 -430 -139 -428
rect -145 -432 -144 -430
rect -142 -432 -139 -430
rect -145 -434 -139 -432
rect -135 -430 -131 -425
rect -135 -432 -134 -430
rect -132 -432 -131 -430
rect -135 -434 -131 -432
rect -233 -447 -211 -446
rect -242 -450 -238 -448
rect -233 -449 -231 -447
rect -229 -448 -211 -447
rect -209 -448 -208 -446
rect -229 -449 -208 -448
rect -203 -446 -193 -445
rect -203 -448 -201 -446
rect -199 -448 -193 -446
rect -203 -449 -193 -448
rect -143 -437 -139 -434
rect -143 -441 -123 -437
rect -127 -445 -123 -441
rect -92 -436 -88 -425
rect -85 -427 -81 -417
rect -85 -429 -84 -427
rect -82 -429 -81 -427
rect -85 -431 -81 -429
rect -92 -437 -74 -436
rect -112 -439 -108 -437
rect -92 -438 -78 -437
rect -112 -441 -111 -439
rect -109 -441 -108 -439
rect -127 -446 -117 -445
rect -127 -448 -121 -446
rect -119 -448 -117 -446
rect -127 -449 -117 -448
rect -112 -446 -108 -441
rect -103 -439 -78 -438
rect -76 -439 -74 -437
rect -103 -441 -101 -439
rect -99 -440 -74 -439
rect -99 -441 -88 -440
rect -103 -442 -88 -441
rect -112 -448 -111 -446
rect -109 -447 -87 -446
rect -109 -448 -91 -447
rect -112 -449 -91 -448
rect -89 -449 -87 -447
rect -233 -450 -208 -449
rect -112 -450 -87 -449
rect -82 -450 -78 -448
rect -242 -452 -241 -450
rect -239 -452 -238 -450
rect -82 -452 -81 -450
rect -79 -452 -78 -450
rect -242 -455 -238 -452
rect -186 -453 -180 -452
rect -186 -455 -184 -453
rect -182 -455 -180 -453
rect -140 -453 -134 -452
rect -140 -455 -138 -453
rect -136 -455 -134 -453
rect -82 -455 -78 -452
rect 420 -359 424 -348
rect 463 -353 467 -348
rect 463 -355 464 -353
rect 466 -355 467 -353
rect 463 -357 467 -355
rect 471 -351 475 -340
rect 471 -353 477 -351
rect 471 -355 474 -353
rect 476 -355 477 -353
rect 471 -357 477 -355
rect 406 -360 424 -359
rect 406 -362 408 -360
rect 410 -361 424 -360
rect 410 -362 435 -361
rect 406 -363 431 -362
rect 420 -364 431 -363
rect 433 -364 435 -362
rect 420 -365 435 -364
rect 440 -362 444 -360
rect 440 -364 441 -362
rect 443 -364 444 -362
rect 440 -369 444 -364
rect 471 -360 475 -357
rect 455 -364 475 -360
rect 455 -368 459 -364
rect 522 -336 526 -332
rect 545 -336 569 -332
rect 509 -337 549 -336
rect 509 -339 523 -337
rect 525 -339 549 -337
rect 509 -340 549 -339
rect 509 -351 513 -340
rect 557 -341 561 -339
rect 565 -340 571 -336
rect 557 -343 558 -341
rect 560 -343 561 -341
rect 557 -344 561 -343
rect 557 -348 564 -344
rect 507 -353 513 -351
rect 507 -355 508 -353
rect 510 -355 513 -353
rect 507 -357 513 -355
rect 517 -353 521 -348
rect 517 -355 518 -353
rect 520 -355 521 -353
rect 517 -357 521 -355
rect 419 -370 441 -369
rect 410 -373 414 -371
rect 419 -372 421 -370
rect 423 -371 441 -370
rect 443 -371 444 -369
rect 423 -372 444 -371
rect 449 -369 459 -368
rect 449 -371 451 -369
rect 453 -371 459 -369
rect 449 -372 459 -371
rect 509 -360 513 -357
rect 509 -364 529 -360
rect 525 -368 529 -364
rect 560 -359 564 -348
rect 567 -350 571 -340
rect 567 -352 568 -350
rect 570 -352 571 -350
rect 567 -354 571 -352
rect 560 -360 578 -359
rect 540 -362 544 -360
rect 560 -361 574 -360
rect 540 -364 541 -362
rect 543 -364 544 -362
rect 525 -369 535 -368
rect 525 -371 531 -369
rect 533 -371 535 -369
rect 525 -372 535 -371
rect 540 -369 544 -364
rect 549 -362 574 -361
rect 576 -362 578 -360
rect 549 -364 551 -362
rect 553 -363 578 -362
rect 553 -364 564 -363
rect 549 -365 564 -364
rect 540 -371 541 -369
rect 543 -370 565 -369
rect 543 -371 561 -370
rect 540 -372 561 -371
rect 563 -372 565 -370
rect 419 -373 444 -372
rect 540 -373 565 -372
rect 570 -373 574 -371
rect 410 -375 411 -373
rect 413 -375 414 -373
rect 570 -375 571 -373
rect 573 -375 574 -373
rect 410 -378 414 -375
rect 466 -376 472 -375
rect 466 -378 468 -376
rect 470 -378 472 -376
rect 512 -376 518 -375
rect 512 -378 514 -376
rect 516 -378 518 -376
rect 570 -378 574 -375
rect 29 -479 31 -477
rect 33 -479 35 -477
rect 29 -484 35 -479
rect 51 -479 53 -477
rect 55 -479 57 -477
rect 29 -486 31 -484
rect 33 -486 35 -484
rect 29 -487 35 -486
rect 40 -485 44 -483
rect 40 -487 41 -485
rect 43 -487 44 -485
rect 51 -484 57 -479
rect 86 -479 88 -477
rect 90 -479 92 -477
rect 86 -480 92 -479
rect 125 -479 127 -477
rect 129 -479 131 -477
rect 125 -480 131 -479
rect 158 -479 160 -477
rect 162 -479 164 -477
rect 51 -486 53 -484
rect 55 -486 57 -484
rect 51 -487 57 -486
rect 107 -484 127 -483
rect 107 -486 109 -484
rect 111 -486 127 -484
rect 107 -487 127 -486
rect 40 -491 44 -487
rect 63 -491 87 -487
rect 27 -492 67 -491
rect 27 -494 41 -492
rect 43 -494 67 -492
rect 27 -495 67 -494
rect 27 -506 31 -495
rect 75 -496 79 -494
rect 83 -495 89 -491
rect 75 -498 76 -496
rect 78 -498 79 -496
rect 75 -499 79 -498
rect 75 -503 82 -499
rect 25 -508 31 -506
rect 25 -510 26 -508
rect 28 -510 31 -508
rect 25 -512 31 -510
rect 35 -508 39 -503
rect 35 -510 36 -508
rect 38 -510 39 -508
rect 35 -512 39 -510
rect 27 -515 31 -512
rect 27 -519 47 -515
rect 43 -523 47 -519
rect 43 -524 51 -523
rect 43 -526 49 -524
rect 43 -527 51 -526
rect 30 -531 36 -530
rect 30 -533 32 -531
rect 34 -533 36 -531
rect 78 -514 82 -503
rect 85 -505 89 -495
rect 85 -507 86 -505
rect 88 -507 89 -505
rect 85 -509 89 -507
rect 78 -515 96 -514
rect 58 -517 62 -515
rect 78 -516 92 -515
rect 58 -519 59 -517
rect 61 -519 62 -517
rect 58 -524 62 -519
rect 67 -517 92 -516
rect 94 -517 96 -515
rect 67 -519 69 -517
rect 71 -518 96 -517
rect 71 -519 82 -518
rect 67 -520 82 -519
rect 123 -491 127 -487
rect 138 -490 139 -487
rect 158 -484 164 -479
rect 180 -479 182 -477
rect 184 -479 186 -477
rect 158 -486 160 -484
rect 162 -486 164 -484
rect 158 -487 164 -486
rect 169 -485 173 -483
rect 169 -487 170 -485
rect 172 -487 173 -485
rect 180 -484 186 -479
rect 215 -479 217 -477
rect 219 -479 221 -477
rect 215 -480 221 -479
rect 249 -479 251 -477
rect 253 -479 255 -477
rect 249 -480 255 -479
rect 284 -479 286 -477
rect 288 -479 290 -477
rect 180 -486 182 -484
rect 184 -486 186 -484
rect 180 -487 186 -486
rect 123 -495 135 -491
rect 131 -507 135 -495
rect 131 -509 132 -507
rect 134 -509 135 -507
rect 131 -514 135 -509
rect 118 -518 135 -514
rect 58 -526 59 -524
rect 61 -525 83 -524
rect 61 -526 79 -525
rect 58 -527 79 -526
rect 81 -527 83 -525
rect 58 -528 83 -527
rect 88 -528 92 -526
rect 107 -522 113 -521
rect 107 -524 109 -522
rect 111 -524 113 -522
rect 88 -530 89 -528
rect 91 -530 92 -528
rect 88 -533 92 -530
rect 107 -533 113 -524
rect 118 -522 122 -518
rect 118 -524 119 -522
rect 121 -524 122 -522
rect 118 -526 122 -524
rect 127 -522 133 -521
rect 127 -524 129 -522
rect 131 -524 133 -522
rect 127 -533 133 -524
rect 169 -491 173 -487
rect 192 -491 216 -487
rect 156 -492 196 -491
rect 156 -494 170 -492
rect 172 -494 196 -492
rect 156 -495 196 -494
rect 156 -506 160 -495
rect 204 -496 208 -494
rect 212 -495 218 -491
rect 204 -498 205 -496
rect 207 -498 208 -496
rect 204 -499 208 -498
rect 204 -503 211 -499
rect 154 -508 160 -506
rect 154 -510 155 -508
rect 157 -510 160 -508
rect 154 -512 160 -510
rect 164 -508 168 -503
rect 164 -510 165 -508
rect 167 -510 168 -508
rect 164 -512 168 -510
rect 156 -515 160 -512
rect 156 -519 176 -515
rect 172 -523 176 -519
rect 207 -514 211 -503
rect 214 -505 218 -495
rect 214 -507 215 -505
rect 217 -507 218 -505
rect 214 -509 218 -507
rect 207 -515 225 -514
rect 187 -517 191 -515
rect 207 -516 221 -515
rect 187 -519 188 -517
rect 190 -519 191 -517
rect 172 -524 182 -523
rect 172 -526 178 -524
rect 180 -526 182 -524
rect 172 -527 182 -526
rect 187 -524 191 -519
rect 196 -517 221 -516
rect 223 -517 225 -515
rect 196 -519 198 -517
rect 200 -518 225 -517
rect 200 -519 211 -518
rect 196 -520 211 -519
rect 187 -526 188 -524
rect 190 -525 212 -524
rect 190 -526 208 -525
rect 187 -527 208 -526
rect 210 -527 212 -525
rect 187 -528 212 -527
rect 217 -528 221 -526
rect 284 -484 290 -479
rect 306 -479 308 -477
rect 310 -479 312 -477
rect 284 -486 286 -484
rect 288 -486 290 -484
rect 284 -487 290 -486
rect 297 -485 301 -483
rect 297 -487 298 -485
rect 300 -487 301 -485
rect 306 -484 312 -479
rect 339 -479 341 -477
rect 343 -479 345 -477
rect 339 -480 345 -479
rect 378 -479 380 -477
rect 382 -479 384 -477
rect 378 -480 384 -479
rect 413 -479 415 -477
rect 417 -479 419 -477
rect 306 -486 308 -484
rect 310 -486 312 -484
rect 306 -487 312 -486
rect 254 -491 278 -487
rect 297 -491 301 -487
rect 343 -484 363 -483
rect 343 -486 359 -484
rect 361 -486 363 -484
rect 343 -487 363 -486
rect 413 -484 419 -479
rect 435 -479 437 -477
rect 439 -479 441 -477
rect 413 -486 415 -484
rect 417 -486 419 -484
rect 413 -487 419 -486
rect 426 -485 430 -483
rect 426 -487 427 -485
rect 429 -487 430 -485
rect 435 -484 441 -479
rect 435 -486 437 -484
rect 439 -486 441 -484
rect 435 -487 441 -486
rect 467 -479 469 -477
rect 471 -479 473 -477
rect 467 -484 473 -479
rect 489 -479 491 -477
rect 493 -479 495 -477
rect 467 -486 469 -484
rect 471 -486 473 -484
rect 467 -487 473 -486
rect 478 -485 482 -483
rect 478 -487 479 -485
rect 481 -487 482 -485
rect 489 -484 495 -479
rect 524 -479 526 -477
rect 528 -479 530 -477
rect 524 -480 530 -479
rect 563 -479 565 -477
rect 567 -479 569 -477
rect 563 -480 569 -479
rect 596 -479 598 -477
rect 600 -479 602 -477
rect 489 -486 491 -484
rect 493 -486 495 -484
rect 489 -487 495 -486
rect 545 -484 565 -483
rect 545 -486 547 -484
rect 549 -486 565 -484
rect 545 -487 565 -486
rect 252 -495 258 -491
rect 274 -492 314 -491
rect 274 -494 298 -492
rect 300 -494 314 -492
rect 252 -505 256 -495
rect 262 -496 266 -494
rect 274 -495 314 -494
rect 262 -498 263 -496
rect 265 -498 266 -496
rect 262 -499 266 -498
rect 252 -507 253 -505
rect 255 -507 256 -505
rect 252 -509 256 -507
rect 259 -503 266 -499
rect 259 -514 263 -503
rect 302 -508 306 -503
rect 302 -510 303 -508
rect 305 -510 306 -508
rect 245 -515 263 -514
rect 245 -517 247 -515
rect 249 -516 263 -515
rect 249 -517 274 -516
rect 245 -518 270 -517
rect 259 -519 270 -518
rect 272 -519 274 -517
rect 259 -520 274 -519
rect 279 -517 283 -515
rect 279 -519 280 -517
rect 282 -519 283 -517
rect 279 -524 283 -519
rect 302 -512 306 -510
rect 310 -506 314 -495
rect 310 -508 316 -506
rect 310 -510 313 -508
rect 315 -510 316 -508
rect 310 -512 316 -510
rect 310 -515 314 -512
rect 294 -519 314 -515
rect 294 -523 298 -519
rect 258 -525 280 -524
rect 249 -528 253 -526
rect 258 -527 260 -525
rect 262 -526 280 -525
rect 282 -526 283 -524
rect 262 -527 283 -526
rect 288 -524 298 -523
rect 288 -526 290 -524
rect 292 -526 298 -524
rect 288 -527 298 -526
rect 331 -490 332 -487
rect 343 -491 347 -487
rect 335 -495 347 -491
rect 335 -507 339 -495
rect 383 -491 407 -487
rect 426 -491 430 -487
rect 335 -509 336 -507
rect 338 -509 339 -507
rect 335 -514 339 -509
rect 381 -495 387 -491
rect 403 -492 443 -491
rect 403 -494 427 -492
rect 429 -494 443 -492
rect 381 -505 385 -495
rect 391 -496 395 -494
rect 403 -495 443 -494
rect 391 -498 392 -496
rect 394 -498 395 -496
rect 391 -499 395 -498
rect 381 -507 382 -505
rect 384 -507 385 -505
rect 381 -509 385 -507
rect 388 -503 395 -499
rect 335 -518 352 -514
rect 258 -528 283 -527
rect 337 -522 343 -521
rect 337 -524 339 -522
rect 341 -524 343 -522
rect 217 -530 218 -528
rect 220 -530 221 -528
rect 159 -531 165 -530
rect 159 -533 161 -531
rect 163 -533 165 -531
rect 217 -533 221 -530
rect 249 -530 250 -528
rect 252 -530 253 -528
rect 249 -533 253 -530
rect 305 -531 311 -530
rect 305 -533 307 -531
rect 309 -533 311 -531
rect 337 -533 343 -524
rect 348 -522 352 -518
rect 348 -524 349 -522
rect 351 -524 352 -522
rect 348 -526 352 -524
rect 357 -522 363 -521
rect 357 -524 359 -522
rect 361 -524 363 -522
rect 357 -533 363 -524
rect 388 -514 392 -503
rect 431 -508 435 -503
rect 431 -510 432 -508
rect 434 -510 435 -508
rect 374 -515 392 -514
rect 374 -517 376 -515
rect 378 -516 392 -515
rect 378 -517 403 -516
rect 374 -518 399 -517
rect 388 -519 399 -518
rect 401 -519 403 -517
rect 388 -520 403 -519
rect 408 -517 412 -515
rect 408 -519 409 -517
rect 411 -519 412 -517
rect 408 -524 412 -519
rect 431 -512 435 -510
rect 439 -506 443 -495
rect 439 -508 445 -506
rect 439 -510 442 -508
rect 444 -510 445 -508
rect 439 -512 445 -510
rect 439 -515 443 -512
rect 423 -519 443 -515
rect 423 -523 427 -519
rect 387 -525 409 -524
rect 378 -528 382 -526
rect 387 -527 389 -525
rect 391 -526 409 -525
rect 411 -526 412 -524
rect 391 -527 412 -526
rect 417 -524 427 -523
rect 417 -526 419 -524
rect 421 -526 427 -524
rect 417 -527 427 -526
rect 478 -491 482 -487
rect 501 -491 525 -487
rect 465 -492 505 -491
rect 465 -494 479 -492
rect 481 -494 505 -492
rect 465 -495 505 -494
rect 465 -506 469 -495
rect 513 -496 517 -494
rect 521 -495 527 -491
rect 513 -498 514 -496
rect 516 -498 517 -496
rect 513 -499 517 -498
rect 513 -503 520 -499
rect 463 -508 469 -506
rect 463 -510 464 -508
rect 466 -510 469 -508
rect 463 -512 469 -510
rect 473 -508 477 -503
rect 473 -510 474 -508
rect 476 -510 477 -508
rect 473 -512 477 -510
rect 465 -515 469 -512
rect 465 -519 485 -515
rect 481 -523 485 -519
rect 516 -514 520 -503
rect 523 -505 527 -495
rect 523 -507 524 -505
rect 526 -507 527 -505
rect 523 -509 527 -507
rect 516 -515 534 -514
rect 496 -517 500 -515
rect 516 -516 530 -515
rect 496 -519 497 -517
rect 499 -519 500 -517
rect 481 -524 491 -523
rect 481 -526 487 -524
rect 489 -526 491 -524
rect 481 -527 491 -526
rect 496 -524 500 -519
rect 505 -517 530 -516
rect 532 -517 534 -515
rect 505 -519 507 -517
rect 509 -518 534 -517
rect 509 -519 520 -518
rect 505 -520 520 -519
rect 561 -491 565 -487
rect 576 -490 577 -487
rect 596 -484 602 -479
rect 618 -479 620 -477
rect 622 -479 624 -477
rect 596 -486 598 -484
rect 600 -486 602 -484
rect 596 -487 602 -486
rect 607 -485 611 -483
rect 607 -487 608 -485
rect 610 -487 611 -485
rect 618 -484 624 -479
rect 653 -479 655 -477
rect 657 -479 659 -477
rect 653 -480 659 -479
rect 688 -479 690 -477
rect 692 -479 694 -477
rect 618 -486 620 -484
rect 622 -486 624 -484
rect 618 -487 624 -486
rect 688 -484 694 -479
rect 710 -479 712 -477
rect 714 -479 716 -477
rect 688 -486 690 -484
rect 692 -486 694 -484
rect 688 -487 694 -486
rect 699 -485 703 -483
rect 699 -487 700 -485
rect 702 -487 703 -485
rect 710 -484 716 -479
rect 745 -479 747 -477
rect 749 -479 751 -477
rect 745 -480 751 -479
rect 710 -486 712 -484
rect 714 -486 716 -484
rect 710 -487 716 -486
rect 561 -495 573 -491
rect 569 -507 573 -495
rect 569 -509 570 -507
rect 572 -509 573 -507
rect 569 -514 573 -509
rect 556 -518 573 -514
rect 496 -526 497 -524
rect 499 -525 521 -524
rect 499 -526 517 -525
rect 496 -527 517 -526
rect 519 -527 521 -525
rect 387 -528 412 -527
rect 496 -528 521 -527
rect 526 -528 530 -526
rect 545 -522 551 -521
rect 545 -524 547 -522
rect 549 -524 551 -522
rect 378 -530 379 -528
rect 381 -530 382 -528
rect 526 -530 527 -528
rect 529 -530 530 -528
rect 378 -533 382 -530
rect 434 -531 440 -530
rect 434 -533 436 -531
rect 438 -533 440 -531
rect 468 -531 474 -530
rect 468 -533 470 -531
rect 472 -533 474 -531
rect 526 -533 530 -530
rect 545 -533 551 -524
rect 556 -522 560 -518
rect 556 -524 557 -522
rect 559 -524 560 -522
rect 556 -526 560 -524
rect 565 -522 571 -521
rect 565 -524 567 -522
rect 569 -524 571 -522
rect 565 -533 571 -524
rect 607 -491 611 -487
rect 630 -491 654 -487
rect 594 -492 634 -491
rect 594 -494 608 -492
rect 610 -494 634 -492
rect 594 -495 634 -494
rect 594 -506 598 -495
rect 642 -496 646 -494
rect 650 -495 656 -491
rect 642 -498 643 -496
rect 645 -498 646 -496
rect 642 -499 646 -498
rect 642 -503 649 -499
rect 592 -508 598 -506
rect 592 -510 593 -508
rect 595 -510 598 -508
rect 592 -512 598 -510
rect 602 -508 606 -503
rect 602 -510 603 -508
rect 605 -510 606 -508
rect 602 -512 606 -510
rect 594 -515 598 -512
rect 594 -519 614 -515
rect 610 -523 614 -519
rect 645 -514 649 -503
rect 652 -505 656 -495
rect 652 -507 653 -505
rect 655 -507 656 -505
rect 652 -509 656 -507
rect 645 -515 663 -514
rect 625 -517 629 -515
rect 645 -516 659 -515
rect 625 -519 626 -517
rect 628 -519 629 -517
rect 610 -524 620 -523
rect 610 -526 616 -524
rect 618 -526 620 -524
rect 610 -527 620 -526
rect 625 -524 629 -519
rect 634 -517 659 -516
rect 661 -517 663 -515
rect 634 -519 636 -517
rect 638 -518 663 -517
rect 638 -519 649 -518
rect 634 -520 649 -519
rect 625 -526 626 -524
rect 628 -525 650 -524
rect 628 -526 646 -525
rect 625 -527 646 -526
rect 648 -527 650 -525
rect 625 -528 650 -527
rect 655 -528 659 -526
rect 699 -491 703 -487
rect 722 -491 746 -487
rect 686 -492 726 -491
rect 686 -494 700 -492
rect 702 -494 726 -492
rect 686 -495 726 -494
rect 686 -506 690 -495
rect 734 -496 738 -494
rect 742 -495 748 -491
rect 734 -498 735 -496
rect 737 -498 738 -496
rect 734 -499 738 -498
rect 734 -503 741 -499
rect 684 -508 690 -506
rect 684 -510 685 -508
rect 687 -510 690 -508
rect 684 -512 690 -510
rect 694 -508 698 -503
rect 694 -510 695 -508
rect 697 -510 698 -508
rect 694 -512 698 -510
rect 686 -515 690 -512
rect 686 -519 706 -515
rect 702 -523 706 -519
rect 737 -514 741 -503
rect 744 -505 748 -495
rect 744 -507 745 -505
rect 747 -507 748 -505
rect 744 -509 748 -507
rect 737 -515 755 -514
rect 717 -517 721 -515
rect 737 -516 751 -515
rect 717 -519 718 -517
rect 720 -519 721 -517
rect 702 -524 712 -523
rect 702 -526 708 -524
rect 710 -526 712 -524
rect 702 -527 712 -526
rect 717 -524 721 -519
rect 726 -517 751 -516
rect 753 -517 755 -515
rect 726 -519 728 -517
rect 730 -518 755 -517
rect 730 -519 741 -518
rect 726 -520 741 -519
rect 717 -526 718 -524
rect 720 -525 742 -524
rect 720 -526 738 -525
rect 717 -527 738 -526
rect 740 -527 742 -525
rect 717 -528 742 -527
rect 747 -528 751 -526
rect 655 -530 656 -528
rect 658 -530 659 -528
rect 747 -530 748 -528
rect 750 -530 751 -528
rect 597 -531 603 -530
rect 597 -533 599 -531
rect 601 -533 603 -531
rect 655 -533 659 -530
rect 689 -531 695 -530
rect 689 -533 691 -531
rect 693 -533 695 -531
rect 747 -533 751 -530
rect -238 -613 -236 -611
rect -234 -613 -232 -611
rect -238 -618 -232 -613
rect -216 -613 -214 -611
rect -212 -613 -210 -611
rect -238 -620 -236 -618
rect -234 -620 -232 -618
rect -238 -621 -232 -620
rect -227 -619 -223 -617
rect -227 -621 -226 -619
rect -224 -621 -223 -619
rect -216 -618 -210 -613
rect -181 -613 -179 -611
rect -177 -613 -175 -611
rect -181 -614 -175 -613
rect -142 -613 -140 -611
rect -138 -613 -136 -611
rect -142 -614 -136 -613
rect -109 -613 -107 -611
rect -105 -613 -103 -611
rect -216 -620 -214 -618
rect -212 -620 -210 -618
rect -216 -621 -210 -620
rect -160 -618 -140 -617
rect -160 -620 -158 -618
rect -156 -620 -140 -618
rect -160 -621 -140 -620
rect -227 -625 -223 -621
rect -204 -625 -180 -621
rect -240 -626 -200 -625
rect -240 -628 -226 -626
rect -224 -628 -200 -626
rect -240 -629 -200 -628
rect -240 -640 -236 -629
rect -192 -630 -188 -628
rect -184 -629 -178 -625
rect -192 -632 -191 -630
rect -189 -632 -188 -630
rect -192 -633 -188 -632
rect -192 -637 -185 -633
rect -242 -642 -236 -640
rect -242 -644 -241 -642
rect -239 -644 -236 -642
rect -242 -646 -236 -644
rect -232 -642 -228 -637
rect -232 -644 -231 -642
rect -229 -644 -228 -642
rect -232 -646 -228 -644
rect -240 -649 -236 -646
rect -240 -653 -220 -649
rect -224 -657 -220 -653
rect -189 -648 -185 -637
rect -182 -639 -178 -629
rect -182 -641 -181 -639
rect -179 -641 -178 -639
rect -182 -643 -178 -641
rect -189 -649 -171 -648
rect -209 -651 -205 -649
rect -189 -650 -175 -649
rect -209 -653 -208 -651
rect -206 -653 -205 -651
rect -224 -658 -214 -657
rect -224 -660 -218 -658
rect -216 -660 -214 -658
rect -224 -661 -214 -660
rect -209 -658 -205 -653
rect -200 -651 -175 -650
rect -173 -651 -171 -649
rect -200 -653 -198 -651
rect -196 -652 -171 -651
rect -196 -653 -185 -652
rect -200 -654 -185 -653
rect -144 -625 -140 -621
rect -129 -624 -128 -621
rect -109 -618 -103 -613
rect -87 -613 -85 -611
rect -83 -613 -81 -611
rect -109 -620 -107 -618
rect -105 -620 -103 -618
rect -109 -621 -103 -620
rect -98 -619 -94 -617
rect -98 -621 -97 -619
rect -95 -621 -94 -619
rect -87 -618 -81 -613
rect -52 -613 -50 -611
rect -48 -613 -46 -611
rect -52 -614 -46 -613
rect -18 -613 -16 -611
rect -14 -613 -12 -611
rect -18 -614 -12 -613
rect 17 -613 19 -611
rect 21 -613 23 -611
rect -87 -620 -85 -618
rect -83 -620 -81 -618
rect -87 -621 -81 -620
rect -144 -629 -132 -625
rect -136 -641 -132 -629
rect -136 -643 -135 -641
rect -133 -643 -132 -641
rect -136 -648 -132 -643
rect -149 -652 -132 -648
rect -209 -660 -208 -658
rect -206 -659 -184 -658
rect -206 -660 -188 -659
rect -209 -661 -188 -660
rect -186 -661 -184 -659
rect -209 -662 -184 -661
rect -179 -662 -175 -660
rect -160 -656 -154 -655
rect -160 -658 -158 -656
rect -156 -658 -154 -656
rect -179 -664 -178 -662
rect -176 -664 -175 -662
rect -237 -665 -231 -664
rect -237 -667 -235 -665
rect -233 -667 -231 -665
rect -179 -667 -175 -664
rect -160 -667 -154 -658
rect -149 -656 -145 -652
rect -149 -658 -148 -656
rect -146 -658 -145 -656
rect -149 -660 -145 -658
rect -140 -656 -134 -655
rect -140 -658 -138 -656
rect -136 -658 -134 -656
rect -140 -667 -134 -658
rect -98 -625 -94 -621
rect -75 -625 -51 -621
rect -111 -626 -71 -625
rect -111 -628 -97 -626
rect -95 -628 -71 -626
rect -111 -629 -71 -628
rect -111 -640 -107 -629
rect -63 -630 -59 -628
rect -55 -629 -49 -625
rect -63 -632 -62 -630
rect -60 -632 -59 -630
rect -63 -633 -59 -632
rect -63 -637 -56 -633
rect -113 -642 -107 -640
rect -113 -644 -112 -642
rect -110 -644 -107 -642
rect -113 -646 -107 -644
rect -103 -642 -99 -637
rect -103 -644 -102 -642
rect -100 -644 -99 -642
rect -103 -646 -99 -644
rect -111 -649 -107 -646
rect -111 -653 -91 -649
rect -95 -657 -91 -653
rect -60 -648 -56 -637
rect -53 -639 -49 -629
rect -53 -641 -52 -639
rect -50 -641 -49 -639
rect -53 -643 -49 -641
rect -60 -649 -42 -648
rect -80 -651 -76 -649
rect -60 -650 -46 -649
rect -80 -653 -79 -651
rect -77 -653 -76 -651
rect -95 -658 -85 -657
rect -95 -660 -89 -658
rect -87 -660 -85 -658
rect -95 -661 -85 -660
rect -80 -658 -76 -653
rect -71 -651 -46 -650
rect -44 -651 -42 -649
rect -71 -653 -69 -651
rect -67 -652 -42 -651
rect -67 -653 -56 -652
rect -71 -654 -56 -653
rect -80 -660 -79 -658
rect -77 -659 -55 -658
rect -77 -660 -59 -659
rect -80 -661 -59 -660
rect -57 -661 -55 -659
rect -80 -662 -55 -661
rect -50 -662 -46 -660
rect 17 -618 23 -613
rect 39 -613 41 -611
rect 43 -613 45 -611
rect 17 -620 19 -618
rect 21 -620 23 -618
rect 17 -621 23 -620
rect 30 -619 34 -617
rect 30 -621 31 -619
rect 33 -621 34 -619
rect 39 -618 45 -613
rect 72 -613 74 -611
rect 76 -613 78 -611
rect 72 -614 78 -613
rect 111 -613 113 -611
rect 115 -613 117 -611
rect 111 -614 117 -613
rect 146 -613 148 -611
rect 150 -613 152 -611
rect 39 -620 41 -618
rect 43 -620 45 -618
rect 39 -621 45 -620
rect -13 -625 11 -621
rect 30 -625 34 -621
rect 76 -618 96 -617
rect 76 -620 92 -618
rect 94 -620 96 -618
rect 76 -621 96 -620
rect 146 -618 152 -613
rect 168 -613 170 -611
rect 172 -613 174 -611
rect 146 -620 148 -618
rect 150 -620 152 -618
rect 146 -621 152 -620
rect 159 -619 163 -617
rect 159 -621 160 -619
rect 162 -621 163 -619
rect 168 -618 174 -613
rect 168 -620 170 -618
rect 172 -620 174 -618
rect 168 -621 174 -620
rect 200 -613 202 -611
rect 204 -613 206 -611
rect 200 -618 206 -613
rect 222 -613 224 -611
rect 226 -613 228 -611
rect 200 -620 202 -618
rect 204 -620 206 -618
rect 200 -621 206 -620
rect 211 -619 215 -617
rect 211 -621 212 -619
rect 214 -621 215 -619
rect 222 -618 228 -613
rect 257 -613 259 -611
rect 261 -613 263 -611
rect 257 -614 263 -613
rect 296 -613 298 -611
rect 300 -613 302 -611
rect 296 -614 302 -613
rect 329 -613 331 -611
rect 333 -613 335 -611
rect 222 -620 224 -618
rect 226 -620 228 -618
rect 222 -621 228 -620
rect 278 -618 298 -617
rect 278 -620 280 -618
rect 282 -620 298 -618
rect 278 -621 298 -620
rect -15 -629 -9 -625
rect 7 -626 47 -625
rect 7 -628 31 -626
rect 33 -628 47 -626
rect -15 -639 -11 -629
rect -5 -630 -1 -628
rect 7 -629 47 -628
rect -5 -632 -4 -630
rect -2 -632 -1 -630
rect -5 -633 -1 -632
rect -15 -641 -14 -639
rect -12 -641 -11 -639
rect -15 -643 -11 -641
rect -8 -637 -1 -633
rect -8 -648 -4 -637
rect 35 -642 39 -637
rect 35 -644 36 -642
rect 38 -644 39 -642
rect -22 -649 -4 -648
rect -22 -651 -20 -649
rect -18 -650 -4 -649
rect -18 -651 7 -650
rect -22 -652 3 -651
rect -8 -653 3 -652
rect 5 -653 7 -651
rect -8 -654 7 -653
rect 12 -651 16 -649
rect 12 -653 13 -651
rect 15 -653 16 -651
rect 12 -658 16 -653
rect 35 -646 39 -644
rect 43 -640 47 -629
rect 43 -642 49 -640
rect 43 -644 46 -642
rect 48 -644 49 -642
rect 43 -646 49 -644
rect 43 -649 47 -646
rect 27 -653 47 -649
rect 27 -657 31 -653
rect -9 -659 13 -658
rect -18 -662 -14 -660
rect -9 -661 -7 -659
rect -5 -660 13 -659
rect 15 -660 16 -658
rect -5 -661 16 -660
rect 21 -658 31 -657
rect 21 -660 23 -658
rect 25 -660 31 -658
rect 21 -661 31 -660
rect 64 -624 65 -621
rect 76 -625 80 -621
rect 68 -629 80 -625
rect 68 -641 72 -629
rect 116 -625 140 -621
rect 159 -625 163 -621
rect 68 -643 69 -641
rect 71 -643 72 -641
rect 68 -648 72 -643
rect 114 -629 120 -625
rect 136 -626 176 -625
rect 136 -628 160 -626
rect 162 -628 176 -626
rect 114 -639 118 -629
rect 124 -630 128 -628
rect 136 -629 176 -628
rect 124 -632 125 -630
rect 127 -632 128 -630
rect 124 -633 128 -632
rect 114 -641 115 -639
rect 117 -641 118 -639
rect 114 -643 118 -641
rect 121 -637 128 -633
rect 68 -652 85 -648
rect -9 -662 16 -661
rect 70 -656 76 -655
rect 70 -658 72 -656
rect 74 -658 76 -656
rect -50 -664 -49 -662
rect -47 -664 -46 -662
rect -108 -665 -102 -664
rect -108 -667 -106 -665
rect -104 -667 -102 -665
rect -50 -667 -46 -664
rect -18 -664 -17 -662
rect -15 -664 -14 -662
rect -18 -667 -14 -664
rect 38 -665 44 -664
rect 38 -667 40 -665
rect 42 -667 44 -665
rect 70 -667 76 -658
rect 81 -656 85 -652
rect 81 -658 82 -656
rect 84 -658 85 -656
rect 81 -660 85 -658
rect 90 -656 96 -655
rect 90 -658 92 -656
rect 94 -658 96 -656
rect 90 -667 96 -658
rect 121 -648 125 -637
rect 164 -642 168 -637
rect 164 -644 165 -642
rect 167 -644 168 -642
rect 107 -649 125 -648
rect 107 -651 109 -649
rect 111 -650 125 -649
rect 111 -651 136 -650
rect 107 -652 132 -651
rect 121 -653 132 -652
rect 134 -653 136 -651
rect 121 -654 136 -653
rect 141 -651 145 -649
rect 141 -653 142 -651
rect 144 -653 145 -651
rect 141 -658 145 -653
rect 164 -646 168 -644
rect 172 -640 176 -629
rect 172 -642 178 -640
rect 172 -644 175 -642
rect 177 -644 178 -642
rect 172 -646 178 -644
rect 172 -649 176 -646
rect 156 -653 176 -649
rect 156 -657 160 -653
rect 120 -659 142 -658
rect 111 -662 115 -660
rect 120 -661 122 -659
rect 124 -660 142 -659
rect 144 -660 145 -658
rect 124 -661 145 -660
rect 150 -658 160 -657
rect 150 -660 152 -658
rect 154 -660 160 -658
rect 150 -661 160 -660
rect 211 -625 215 -621
rect 234 -625 258 -621
rect 198 -626 238 -625
rect 198 -628 212 -626
rect 214 -628 238 -626
rect 198 -629 238 -628
rect 198 -640 202 -629
rect 246 -630 250 -628
rect 254 -629 260 -625
rect 246 -632 247 -630
rect 249 -632 250 -630
rect 246 -633 250 -632
rect 246 -637 253 -633
rect 196 -642 202 -640
rect 196 -644 197 -642
rect 199 -644 202 -642
rect 196 -646 202 -644
rect 206 -642 210 -637
rect 206 -644 207 -642
rect 209 -644 210 -642
rect 206 -646 210 -644
rect 198 -649 202 -646
rect 198 -653 218 -649
rect 214 -657 218 -653
rect 249 -648 253 -637
rect 256 -639 260 -629
rect 256 -641 257 -639
rect 259 -641 260 -639
rect 256 -643 260 -641
rect 249 -649 267 -648
rect 229 -651 233 -649
rect 249 -650 263 -649
rect 229 -653 230 -651
rect 232 -653 233 -651
rect 214 -658 224 -657
rect 214 -660 220 -658
rect 222 -660 224 -658
rect 214 -661 224 -660
rect 229 -658 233 -653
rect 238 -651 263 -650
rect 265 -651 267 -649
rect 238 -653 240 -651
rect 242 -652 267 -651
rect 242 -653 253 -652
rect 238 -654 253 -653
rect 294 -625 298 -621
rect 309 -624 310 -621
rect 329 -618 335 -613
rect 351 -613 353 -611
rect 355 -613 357 -611
rect 329 -620 331 -618
rect 333 -620 335 -618
rect 329 -621 335 -620
rect 340 -619 344 -617
rect 340 -621 341 -619
rect 343 -621 344 -619
rect 351 -618 357 -613
rect 386 -613 388 -611
rect 390 -613 392 -611
rect 386 -614 392 -613
rect 421 -613 423 -611
rect 425 -613 427 -611
rect 351 -620 353 -618
rect 355 -620 357 -618
rect 351 -621 357 -620
rect 421 -618 427 -613
rect 443 -613 445 -611
rect 447 -613 449 -611
rect 421 -620 423 -618
rect 425 -620 427 -618
rect 421 -621 427 -620
rect 432 -619 436 -617
rect 432 -621 433 -619
rect 435 -621 436 -619
rect 443 -618 449 -613
rect 478 -613 480 -611
rect 482 -613 484 -611
rect 478 -614 484 -613
rect 443 -620 445 -618
rect 447 -620 449 -618
rect 443 -621 449 -620
rect 294 -629 306 -625
rect 302 -641 306 -629
rect 302 -643 303 -641
rect 305 -643 306 -641
rect 302 -648 306 -643
rect 289 -652 306 -648
rect 229 -660 230 -658
rect 232 -659 254 -658
rect 232 -660 250 -659
rect 229 -661 250 -660
rect 252 -661 254 -659
rect 120 -662 145 -661
rect 229 -662 254 -661
rect 259 -662 263 -660
rect 278 -656 284 -655
rect 278 -658 280 -656
rect 282 -658 284 -656
rect 111 -664 112 -662
rect 114 -664 115 -662
rect 259 -664 260 -662
rect 262 -664 263 -662
rect 111 -667 115 -664
rect 167 -665 173 -664
rect 167 -667 169 -665
rect 171 -667 173 -665
rect 201 -665 207 -664
rect 201 -667 203 -665
rect 205 -667 207 -665
rect 259 -667 263 -664
rect 278 -667 284 -658
rect 289 -656 293 -652
rect 289 -658 290 -656
rect 292 -658 293 -656
rect 289 -660 293 -658
rect 298 -656 304 -655
rect 298 -658 300 -656
rect 302 -658 304 -656
rect 298 -667 304 -658
rect 340 -625 344 -621
rect 363 -625 387 -621
rect 327 -626 367 -625
rect 327 -628 341 -626
rect 343 -628 367 -626
rect 327 -629 367 -628
rect 327 -640 331 -629
rect 375 -630 379 -628
rect 383 -629 389 -625
rect 375 -632 376 -630
rect 378 -632 379 -630
rect 375 -633 379 -632
rect 375 -637 382 -633
rect 325 -642 331 -640
rect 325 -644 326 -642
rect 328 -644 331 -642
rect 325 -646 331 -644
rect 335 -642 339 -637
rect 335 -644 336 -642
rect 338 -644 339 -642
rect 335 -646 339 -644
rect 327 -649 331 -646
rect 327 -653 347 -649
rect 343 -657 347 -653
rect 378 -648 382 -637
rect 385 -639 389 -629
rect 385 -641 386 -639
rect 388 -641 389 -639
rect 385 -643 389 -641
rect 378 -649 396 -648
rect 358 -651 362 -649
rect 378 -650 392 -649
rect 358 -653 359 -651
rect 361 -653 362 -651
rect 343 -658 353 -657
rect 343 -660 349 -658
rect 351 -660 353 -658
rect 343 -661 353 -660
rect 358 -658 362 -653
rect 367 -651 392 -650
rect 394 -651 396 -649
rect 367 -653 369 -651
rect 371 -652 396 -651
rect 371 -653 382 -652
rect 367 -654 382 -653
rect 358 -660 359 -658
rect 361 -659 383 -658
rect 361 -660 379 -659
rect 358 -661 379 -660
rect 381 -661 383 -659
rect 358 -662 383 -661
rect 388 -662 392 -660
rect 432 -625 436 -621
rect 455 -625 479 -621
rect 419 -626 459 -625
rect 419 -628 433 -626
rect 435 -628 459 -626
rect 419 -629 459 -628
rect 419 -640 423 -629
rect 467 -630 471 -628
rect 475 -629 481 -625
rect 467 -632 468 -630
rect 470 -632 471 -630
rect 467 -633 471 -632
rect 467 -637 474 -633
rect 417 -642 423 -640
rect 417 -644 418 -642
rect 420 -644 423 -642
rect 417 -646 423 -644
rect 427 -642 431 -637
rect 427 -644 428 -642
rect 430 -644 431 -642
rect 427 -646 431 -644
rect 419 -649 423 -646
rect 419 -653 439 -649
rect 435 -657 439 -653
rect 470 -648 474 -637
rect 477 -639 481 -629
rect 477 -641 478 -639
rect 480 -641 481 -639
rect 477 -643 481 -641
rect 470 -649 488 -648
rect 450 -651 454 -649
rect 470 -650 484 -649
rect 450 -653 451 -651
rect 453 -653 454 -651
rect 435 -658 445 -657
rect 435 -660 441 -658
rect 443 -660 445 -658
rect 435 -661 445 -660
rect 450 -658 454 -653
rect 459 -651 484 -650
rect 486 -651 488 -649
rect 459 -653 461 -651
rect 463 -652 488 -651
rect 463 -653 474 -652
rect 459 -654 474 -653
rect 450 -660 451 -658
rect 453 -659 475 -658
rect 453 -660 471 -659
rect 450 -661 471 -660
rect 473 -661 475 -659
rect 450 -662 475 -661
rect 480 -662 484 -660
rect 388 -664 389 -662
rect 391 -664 392 -662
rect 480 -664 481 -662
rect 483 -664 484 -662
rect 330 -665 336 -664
rect 330 -667 332 -665
rect 334 -667 336 -665
rect 388 -667 392 -664
rect 422 -665 428 -664
rect 422 -667 424 -665
rect 426 -667 428 -665
rect 480 -667 484 -664
<< via1 >>
rect 268 151 270 153
rect 311 150 313 152
rect 354 150 356 152
rect 415 182 417 184
rect 398 141 400 143
rect 307 70 309 72
rect 315 58 317 60
rect 267 52 269 54
rect 417 70 419 72
rect 368 59 370 61
rect 395 62 397 64
rect 352 50 354 52
rect 449 53 451 55
rect -228 -60 -226 -58
rect -252 -91 -250 -89
rect -209 -92 -207 -90
rect -123 -68 -121 -66
rect -166 -92 -164 -90
rect -99 -59 -97 -57
rect 129 -101 131 -99
rect 19 -116 21 -114
rect 66 -125 68 -123
rect 98 -125 100 -123
rect 50 -134 52 -132
rect 106 -116 108 -114
rect 123 -117 125 -115
rect -213 -172 -211 -170
rect -253 -182 -251 -180
rect -205 -184 -203 -182
rect -103 -172 -101 -170
rect -152 -183 -150 -181
rect -125 -180 -123 -178
rect -168 -196 -166 -194
rect -71 -191 -69 -189
rect 148 -116 150 -114
rect 187 -117 189 -115
rect 179 -134 181 -132
rect 226 -141 228 -139
rect 285 -117 287 -115
rect 316 -116 318 -114
rect 285 -134 287 -132
rect 238 -141 240 -139
rect 326 -109 328 -107
rect 341 -117 343 -115
rect 358 -116 360 -114
rect 366 -125 368 -123
rect 398 -125 400 -123
rect 414 -128 416 -126
rect 445 -116 447 -114
rect 457 -116 459 -114
rect 505 -125 507 -123
rect 488 -129 490 -127
rect 536 -125 538 -123
rect 544 -116 546 -114
rect 561 -117 563 -115
rect 576 -107 578 -105
rect 586 -116 588 -114
rect 623 -117 625 -115
rect 617 -134 619 -132
rect 665 -138 667 -136
rect 692 -117 694 -115
rect 676 -126 678 -124
rect 700 -125 702 -123
rect 757 -126 759 -123
rect 638 -213 640 -211
rect 775 -213 777 -211
rect -251 -343 -249 -341
rect -208 -344 -206 -342
rect -165 -344 -163 -342
rect -104 -312 -102 -310
rect -122 -344 -120 -342
rect 419 -235 421 -233
rect 433 -259 435 -257
rect 401 -266 403 -264
rect 444 -267 446 -265
rect 487 -267 489 -265
rect 554 -235 556 -233
rect 591 -308 593 -306
rect 440 -347 442 -345
rect 400 -358 402 -356
rect -212 -424 -210 -422
rect -252 -434 -250 -432
rect -204 -436 -202 -434
rect -102 -424 -100 -422
rect -151 -435 -149 -433
rect -124 -432 -122 -430
rect -167 -447 -165 -445
rect -70 -435 -68 -433
rect 448 -359 450 -357
rect 550 -347 552 -345
rect 501 -358 503 -356
rect 528 -355 530 -353
rect 484 -371 486 -369
rect 411 -384 413 -382
rect 21 -501 23 -499
rect 68 -510 70 -508
rect 100 -510 102 -508
rect 108 -501 110 -499
rect 125 -502 127 -500
rect 150 -501 152 -499
rect 189 -502 191 -500
rect 181 -519 183 -517
rect 228 -526 230 -524
rect 287 -502 289 -500
rect 318 -501 320 -499
rect 287 -519 289 -517
rect 240 -526 242 -524
rect 328 -494 330 -492
rect 343 -502 345 -500
rect 360 -501 362 -499
rect 368 -510 370 -508
rect 400 -510 402 -508
rect 447 -501 449 -499
rect 416 -518 418 -516
rect 459 -501 461 -499
rect 506 -510 508 -508
rect 538 -510 540 -508
rect 490 -519 492 -517
rect 546 -501 548 -499
rect 563 -502 565 -500
rect 578 -492 580 -490
rect 588 -501 590 -499
rect 625 -502 627 -500
rect 619 -519 621 -517
rect 718 -502 720 -500
rect 678 -511 680 -509
rect 702 -510 704 -508
rect -246 -635 -244 -633
rect -199 -644 -197 -642
rect -167 -644 -165 -642
rect -215 -653 -213 -651
rect -159 -635 -157 -633
rect -142 -636 -140 -634
rect -117 -635 -115 -633
rect -78 -636 -76 -634
rect -86 -653 -84 -651
rect 20 -636 22 -634
rect 51 -635 53 -633
rect 20 -653 22 -651
rect 61 -628 63 -626
rect 76 -636 78 -634
rect 93 -635 95 -633
rect 101 -644 103 -642
rect 129 -644 131 -642
rect 180 -635 182 -633
rect 149 -653 151 -651
rect 192 -635 194 -633
rect 240 -644 242 -642
rect 271 -644 273 -642
rect 223 -653 225 -651
rect 279 -635 281 -633
rect 296 -636 298 -634
rect 311 -626 313 -624
rect 321 -635 323 -633
rect 358 -636 360 -634
rect 352 -653 354 -651
rect 453 -636 455 -634
rect 411 -645 413 -643
rect 445 -644 447 -642
rect 149 -671 151 -669
<< via2 >>
rect -31 197 -29 199
rect 495 53 497 55
rect 253 5 255 7
rect 352 -11 354 -9
rect 688 -12 690 -10
rect 654 -29 656 -27
rect 141 -101 143 -99
rect 285 -109 287 -107
rect 564 -104 566 -102
rect 56 -134 58 -132
rect 227 -167 229 -165
rect 238 -167 240 -165
rect 67 -180 69 -178
rect 406 -128 408 -126
rect 495 -129 497 -127
rect 398 -180 400 -178
rect 725 -13 727 -11
rect 669 -173 671 -170
rect 65 -216 67 -214
rect 692 -236 694 -234
rect 341 -259 343 -257
rect -32 -287 -30 -285
rect -46 -482 -44 -480
rect 411 -400 413 -398
rect 497 -400 499 -398
rect 529 -400 531 -398
rect 422 -412 424 -410
rect 287 -494 289 -492
rect 566 -489 568 -487
rect 68 -521 70 -519
rect 400 -521 402 -519
rect 410 -518 412 -516
rect 497 -519 499 -517
rect 184 -573 186 -571
rect 229 -573 231 -571
rect 506 -523 508 -521
rect 453 -561 455 -559
rect 20 -628 22 -626
rect 299 -623 301 -621
rect -222 -653 -220 -651
rect 217 -648 219 -646
rect 5 -710 7 -708
<< via3 >>
rect 388 4 391 6
rect 495 -40 497 -38
rect 406 -117 408 -115
rect 495 -117 497 -115
rect -47 -526 -45 -524
rect 385 -412 387 -410
rect 497 -418 499 -416
rect 516 -451 518 -449
rect 410 -458 412 -456
rect 410 -504 412 -502
rect 384 -521 386 -519
rect 497 -508 499 -506
rect 515 -524 517 -522
rect 228 -590 230 -588
rect 217 -639 219 -637
rect -47 -710 -45 -708
<< labels >>
rlabel polyct1 -233 -59 -233 -59 1 y1
rlabel polyct1 -104 -59 -104 -59 1 yo
rlabel alu1 51 -128 51 -128 1 a4
rlabel alu1 67 -123 67 -123 1 b4
rlabel alu1 172 -116 172 -116 1 ci4
rlabel alu1 228 -124 228 -124 1 so4
rlabel alu1 238 -124 238 -124 1 so3
rlabel alu1 294 -116 294 -116 1 ci3
rlabel alu1 139 -124 139 -124 1 co4
rlabel alu1 327 -124 327 -124 1 co3
rlabel alu1 577 -124 577 -124 1 co2
rlabel alu1 666 -124 666 -124 1 so2
rlabel alu1 610 -116 610 -116 1 ci2
rlabel via1 489 -128 489 -128 1 a2
rlabel alu1 415 -128 415 -128 1 a3
rlabel via1 399 -124 399 -124 1 b3
rlabel alu1 505 -124 505 -124 1 b2
rlabel via1 758 -124 758 -124 1 so1
rlabel alu2 678 -112 678 -112 1 co1
rlabel alu1 702 -124 702 -124 1 a1
rlabel alu1 694 -116 694 -116 1 b1
rlabel polyct1 -95 -91 -95 -91 1 x2
rlabel polyct1 -224 -91 -224 -91 1 x3
rlabel polyct1 -94 -343 -94 -343 1 x2
rlabel polyct1 -103 -311 -103 -311 1 y2
rlabel polyct1 -232 -311 -232 -311 1 y3
rlabel alu1 583 -354 583 -354 1 m1
rlabel alu1 531 -259 531 -259 1 m0
rlabel alu1 401 -354 401 -354 1 p2
rlabel alu1 481 -342 481 -342 1 p3
rlabel polyct1 558 -266 558 -266 1 xo
rlabel polyct1 549 -234 549 -234 1 yo
rlabel polyct1 429 -266 429 -266 1 x1
rlabel polyct1 296 151 296 151 1 x1
rlabel polyct1 425 151 425 151 1 xo
rlabel polyct1 416 183 416 183 1 y2
rlabel polyct1 287 183 287 183 1 y3
rlabel alu1 760 -509 760 -509 1 m2
rlabel alu1 668 -509 668 -509 1 m3
rlabel via1 69 -508 69 -508 1 b41
rlabel alu1 141 -509 141 -509 1 co41
rlabel alu1 174 -501 174 -501 1 ci41
rlabel alu1 230 -509 230 -509 1 so41
rlabel alu1 240 -509 240 -509 1 so31
rlabel alu1 296 -501 296 -501 1 ci31
rlabel alu1 329 -509 329 -509 1 co31
rlabel via1 401 -509 401 -509 1 b31
rlabel alu1 491 -513 491 -513 1 a21
rlabel via1 507 -509 507 -509 1 b21
rlabel alu1 579 -509 579 -509 1 co21
rlabel alu1 612 -501 612 -501 1 ci21
rlabel alu2 680 -497 680 -497 1 co11
rlabel alu1 696 -501 696 -501 1 b11
rlabel via1 704 -509 704 -509 1 a11
rlabel alu1 268 63 268 63 1 p21
rlabel alu1 348 75 348 75 1 p31
rlabel alu1 450 63 450 63 1 p11
rlabel alu1 -70 -179 -70 -179 1 p13
rlabel alu1 -172 -167 -172 -167 1 p33
rlabel alu2 -252 -179 -252 -179 1 p23
rlabel alu2 -251 -431 -251 -431 1 p22
rlabel alu1 -171 -419 -171 -419 1 p32
rlabel alu2 -69 -431 -69 -431 1 p12
rlabel polyct1 -223 -343 -223 -343 1 x3
rlabel via1 420 -234 420 -234 1 y1
rlabel alu1 332 258 332 258 1 vdd
rlabel alu1 446 -745 446 -745 1 Gnd
rlabel alu1 -81 -607 -81 -607 4 vdd
rlabel alu1 -81 -671 -81 -671 1 Gnd
rlabel alu1 -37 -643 -37 -643 1 m7
rlabel alu1 -27 -643 -27 -643 1 m6
rlabel alu1 -214 -647 -214 -647 1 a42
rlabel poly -192 -648 -192 -648 1 b42
rlabel alu1 29 -635 29 -635 1 ci32
rlabel alu1 134 -643 134 -643 1 b32
rlabel alu1 150 -647 150 -647 1 a32
rlabel alu1 224 -647 224 -647 1 a22
rlabel alu1 240 -643 240 -643 1 b22
rlabel alu1 62 -643 62 -643 1 co32
rlabel alu1 429 -635 429 -635 1 b12
rlabel alu1 437 -643 437 -643 1 a12
rlabel alu2 413 -631 413 -631 1 co12
rlabel alu1 493 -643 493 -643 1 m4
rlabel alu1 401 -643 401 -643 1 m5
rlabel alu1 345 -635 345 -635 1 ci22
rlabel alu1 312 -643 312 -643 1 co22
rlabel alu1 -93 -635 -93 -635 1 ci42
rlabel alu1 -126 -643 -126 -643 1 co42
<< end >>
